magic
tech sky130B
magscale 1 2
timestamp 1662317630
<< locali >>
rect 250740 136740 250860 136760
rect 250740 134420 250760 136740
rect 250840 134420 250860 136740
rect 250740 134400 250860 134420
rect 128660 86660 128700 86840
rect 129200 86660 129240 86840
rect 128660 85060 128700 85220
rect 129200 85060 129240 85220
rect 128520 84970 128550 85060
rect 129330 84970 129360 85060
rect 128520 84960 129360 84970
<< viali >>
rect 250760 134420 250840 136740
rect 128550 84970 129330 85060
<< metal1 >>
rect 250740 136750 250900 136760
rect 250740 136650 250750 136750
rect 250570 136600 250750 136650
rect 250740 136030 250750 136600
rect 250570 135980 250750 136030
rect 250500 135910 250660 135920
rect 250500 135260 250510 135910
rect 250570 135870 250660 135910
rect 250570 135840 250590 135870
rect 250740 135840 250750 135980
rect 250570 135340 250580 135840
rect 250640 135340 250750 135840
rect 250570 135300 250590 135340
rect 250570 135260 250660 135300
rect 250500 135250 250660 135260
rect 250740 135190 250750 135340
rect 250560 135150 250750 135190
rect 250740 134580 250750 135150
rect 250570 134530 250750 134580
rect 250740 134410 250750 134530
rect 250890 134410 250900 136750
rect 250740 134400 250900 134410
rect 233000 123900 235000 124000
rect 233000 123880 233120 123900
rect 233380 123880 233620 123900
rect 233880 123880 234120 123900
rect 234380 123880 234620 123900
rect 234880 123880 235000 123900
rect 233000 123620 233100 123880
rect 233400 123620 233600 123880
rect 233900 123620 234100 123880
rect 234400 123620 234600 123880
rect 234900 123620 235000 123880
rect 233000 123600 233120 123620
rect 233380 123600 233620 123620
rect 233880 123600 234120 123620
rect 234380 123600 234620 123620
rect 234880 123600 235000 123620
rect 233000 123400 235000 123600
rect 233000 123380 233120 123400
rect 233380 123380 233620 123400
rect 233880 123380 234120 123400
rect 234380 123380 234620 123400
rect 234880 123380 235000 123400
rect 233000 123120 233100 123380
rect 233400 123120 233600 123380
rect 233900 123120 234100 123380
rect 234400 123120 234600 123380
rect 234900 123120 235000 123380
rect 233000 123100 233120 123120
rect 233380 123100 233620 123120
rect 233880 123100 234120 123120
rect 234380 123100 234620 123120
rect 234880 123100 235000 123120
rect 233000 122900 235000 123100
rect 233000 122880 233120 122900
rect 233380 122880 233620 122900
rect 233880 122880 234120 122900
rect 234380 122880 234620 122900
rect 234880 122880 235000 122900
rect 233000 122620 233100 122880
rect 233400 122620 233600 122880
rect 233900 122620 234100 122880
rect 234400 122620 234600 122880
rect 234900 122620 235000 122880
rect 233000 122600 233120 122620
rect 233380 122600 233620 122620
rect 233880 122600 234120 122620
rect 234380 122600 234620 122620
rect 234880 122600 235000 122620
rect 233000 122400 235000 122600
rect 233000 122380 233120 122400
rect 233380 122380 233620 122400
rect 233880 122380 234120 122400
rect 234380 122380 234620 122400
rect 234880 122380 235000 122400
rect 233000 122120 233100 122380
rect 233400 122120 233600 122380
rect 233900 122120 234100 122380
rect 234400 122120 234600 122380
rect 234900 122120 235000 122380
rect 233000 122100 233120 122120
rect 233380 122100 233620 122120
rect 233880 122100 234120 122120
rect 234380 122100 234620 122120
rect 234880 122100 235000 122120
rect 233000 122000 235000 122100
rect 14000 121900 58000 122000
rect 14000 121880 14120 121900
rect 14380 121880 14620 121900
rect 14880 121880 15120 121900
rect 15380 121880 15620 121900
rect 15880 121880 16120 121900
rect 16380 121880 16620 121900
rect 16880 121880 17120 121900
rect 17380 121880 17620 121900
rect 17880 121880 18120 121900
rect 18380 121880 18620 121900
rect 18880 121880 19120 121900
rect 19380 121880 19620 121900
rect 19880 121880 20120 121900
rect 20380 121880 20620 121900
rect 20880 121880 21120 121900
rect 21380 121880 21620 121900
rect 21880 121880 22120 121900
rect 22380 121880 22620 121900
rect 22880 121880 23120 121900
rect 23380 121880 23620 121900
rect 23880 121880 24120 121900
rect 24380 121880 24620 121900
rect 24880 121880 25120 121900
rect 25380 121880 25620 121900
rect 25880 121880 26120 121900
rect 26380 121880 26620 121900
rect 26880 121880 27120 121900
rect 27380 121880 27620 121900
rect 27880 121880 28120 121900
rect 28380 121880 28620 121900
rect 28880 121880 29120 121900
rect 29380 121880 29620 121900
rect 29880 121880 30120 121900
rect 30380 121880 30620 121900
rect 30880 121880 31120 121900
rect 31380 121880 31620 121900
rect 31880 121880 32120 121900
rect 32380 121880 32620 121900
rect 32880 121880 33120 121900
rect 33380 121880 33620 121900
rect 33880 121880 34120 121900
rect 34380 121880 34620 121900
rect 34880 121880 35120 121900
rect 35380 121880 35620 121900
rect 35880 121880 36120 121900
rect 36380 121880 36620 121900
rect 36880 121880 37120 121900
rect 37380 121880 37620 121900
rect 37880 121880 38120 121900
rect 38380 121880 38620 121900
rect 38880 121880 39120 121900
rect 39380 121880 39620 121900
rect 39880 121880 40120 121900
rect 40380 121880 40620 121900
rect 40880 121880 41120 121900
rect 41380 121880 41620 121900
rect 41880 121880 42120 121900
rect 42380 121880 42620 121900
rect 42880 121880 43120 121900
rect 43380 121880 43620 121900
rect 43880 121880 44120 121900
rect 44380 121880 44620 121900
rect 44880 121880 45120 121900
rect 45380 121880 45620 121900
rect 45880 121880 46120 121900
rect 46380 121880 46620 121900
rect 46880 121880 47120 121900
rect 47380 121880 47620 121900
rect 47880 121880 48120 121900
rect 48380 121880 48620 121900
rect 48880 121880 49120 121900
rect 49380 121880 49620 121900
rect 49880 121880 50120 121900
rect 50380 121880 50620 121900
rect 50880 121880 51120 121900
rect 51380 121880 51620 121900
rect 51880 121880 52120 121900
rect 52380 121880 52620 121900
rect 52880 121880 53120 121900
rect 53380 121880 53620 121900
rect 53880 121880 54120 121900
rect 54380 121880 54620 121900
rect 54880 121880 55120 121900
rect 55380 121880 55620 121900
rect 55880 121880 56120 121900
rect 56380 121880 56620 121900
rect 56880 121880 57120 121900
rect 57380 121880 57620 121900
rect 57880 121880 58000 121900
rect 14000 121620 14100 121880
rect 14400 121620 14600 121880
rect 14900 121620 15100 121880
rect 15400 121620 15600 121880
rect 15900 121620 16100 121880
rect 16400 121620 16600 121880
rect 16900 121620 17100 121880
rect 17400 121620 17600 121880
rect 17900 121620 18100 121880
rect 18400 121620 18600 121880
rect 18900 121620 19100 121880
rect 19400 121620 19600 121880
rect 19900 121620 20100 121880
rect 20400 121620 20600 121880
rect 20900 121620 21100 121880
rect 21400 121620 21600 121880
rect 21900 121620 22100 121880
rect 22400 121620 22600 121880
rect 22900 121620 23100 121880
rect 23400 121620 23600 121880
rect 23900 121620 24100 121880
rect 24400 121620 24600 121880
rect 24900 121620 25100 121880
rect 25400 121620 25600 121880
rect 25900 121620 26100 121880
rect 26400 121620 26600 121880
rect 26900 121620 27100 121880
rect 27400 121620 27600 121880
rect 27900 121620 28100 121880
rect 28400 121620 28600 121880
rect 28900 121620 29100 121880
rect 29400 121620 29600 121880
rect 29900 121620 30100 121880
rect 30400 121620 30600 121880
rect 30900 121620 31100 121880
rect 31400 121620 31600 121880
rect 31900 121620 32100 121880
rect 32400 121620 32600 121880
rect 32900 121620 33100 121880
rect 33400 121620 33600 121880
rect 33900 121620 34100 121880
rect 34400 121620 34600 121880
rect 34900 121620 35100 121880
rect 35400 121620 35600 121880
rect 35900 121620 36100 121880
rect 36400 121620 36600 121880
rect 36900 121620 37100 121880
rect 37400 121620 37600 121880
rect 37900 121620 38100 121880
rect 38400 121620 38600 121880
rect 38900 121620 39100 121880
rect 39400 121620 39600 121880
rect 39900 121620 40100 121880
rect 40400 121620 40600 121880
rect 40900 121620 41100 121880
rect 41400 121620 41600 121880
rect 41900 121620 42100 121880
rect 42400 121620 42600 121880
rect 42900 121620 43100 121880
rect 43400 121620 43600 121880
rect 43900 121620 44100 121880
rect 44400 121620 44600 121880
rect 44900 121620 45100 121880
rect 45400 121620 45600 121880
rect 45900 121620 46100 121880
rect 46400 121620 46600 121880
rect 46900 121620 47100 121880
rect 47400 121620 47600 121880
rect 47900 121620 48100 121880
rect 48400 121620 48600 121880
rect 48900 121620 49100 121880
rect 49400 121620 49600 121880
rect 49900 121620 50100 121880
rect 50400 121620 50600 121880
rect 50900 121620 51100 121880
rect 51400 121620 51600 121880
rect 51900 121620 52100 121880
rect 52400 121620 52600 121880
rect 52900 121620 53100 121880
rect 53400 121620 53600 121880
rect 53900 121620 54100 121880
rect 54400 121620 54600 121880
rect 54900 121620 55100 121880
rect 55400 121620 55600 121880
rect 55900 121620 56100 121880
rect 56400 121620 56600 121880
rect 56900 121620 57100 121880
rect 57400 121620 57600 121880
rect 57900 121620 58000 121880
rect 14000 121600 14120 121620
rect 14380 121600 14620 121620
rect 14880 121600 15120 121620
rect 15380 121600 15620 121620
rect 15880 121600 16120 121620
rect 16380 121600 16620 121620
rect 16880 121600 17120 121620
rect 17380 121600 17620 121620
rect 17880 121600 18120 121620
rect 18380 121600 18620 121620
rect 18880 121600 19120 121620
rect 19380 121600 19620 121620
rect 19880 121600 20120 121620
rect 20380 121600 20620 121620
rect 20880 121600 21120 121620
rect 21380 121600 21620 121620
rect 21880 121600 22120 121620
rect 22380 121600 22620 121620
rect 22880 121600 23120 121620
rect 23380 121600 23620 121620
rect 23880 121600 24120 121620
rect 24380 121600 24620 121620
rect 24880 121600 25120 121620
rect 25380 121600 25620 121620
rect 25880 121600 26120 121620
rect 26380 121600 26620 121620
rect 26880 121600 27120 121620
rect 27380 121600 27620 121620
rect 27880 121600 28120 121620
rect 28380 121600 28620 121620
rect 28880 121600 29120 121620
rect 29380 121600 29620 121620
rect 29880 121600 30120 121620
rect 30380 121600 30620 121620
rect 30880 121600 31120 121620
rect 31380 121600 31620 121620
rect 31880 121600 32120 121620
rect 32380 121600 32620 121620
rect 32880 121600 33120 121620
rect 33380 121600 33620 121620
rect 33880 121600 34120 121620
rect 34380 121600 34620 121620
rect 34880 121600 35120 121620
rect 35380 121600 35620 121620
rect 35880 121600 36120 121620
rect 36380 121600 36620 121620
rect 36880 121600 37120 121620
rect 37380 121600 37620 121620
rect 37880 121600 38120 121620
rect 38380 121600 38620 121620
rect 38880 121600 39120 121620
rect 39380 121600 39620 121620
rect 39880 121600 40120 121620
rect 40380 121600 40620 121620
rect 40880 121600 41120 121620
rect 41380 121600 41620 121620
rect 41880 121600 42120 121620
rect 42380 121600 42620 121620
rect 42880 121600 43120 121620
rect 43380 121600 43620 121620
rect 43880 121600 44120 121620
rect 44380 121600 44620 121620
rect 44880 121600 45120 121620
rect 45380 121600 45620 121620
rect 45880 121600 46120 121620
rect 46380 121600 46620 121620
rect 46880 121600 47120 121620
rect 47380 121600 47620 121620
rect 47880 121600 48120 121620
rect 48380 121600 48620 121620
rect 48880 121600 49120 121620
rect 49380 121600 49620 121620
rect 49880 121600 50120 121620
rect 50380 121600 50620 121620
rect 50880 121600 51120 121620
rect 51380 121600 51620 121620
rect 51880 121600 52120 121620
rect 52380 121600 52620 121620
rect 52880 121600 53120 121620
rect 53380 121600 53620 121620
rect 53880 121600 54120 121620
rect 54380 121600 54620 121620
rect 54880 121600 55120 121620
rect 55380 121600 55620 121620
rect 55880 121600 56120 121620
rect 56380 121600 56620 121620
rect 56880 121600 57120 121620
rect 57380 121600 57620 121620
rect 57880 121600 58000 121620
rect 14000 121400 58000 121600
rect 14000 121380 14120 121400
rect 14380 121380 14620 121400
rect 14880 121380 15120 121400
rect 15380 121380 15620 121400
rect 15880 121380 16120 121400
rect 16380 121380 16620 121400
rect 16880 121380 17120 121400
rect 17380 121380 17620 121400
rect 17880 121380 18120 121400
rect 18380 121380 18620 121400
rect 18880 121380 19120 121400
rect 19380 121380 19620 121400
rect 19880 121380 20120 121400
rect 20380 121380 20620 121400
rect 20880 121380 21120 121400
rect 21380 121380 21620 121400
rect 21880 121380 22120 121400
rect 22380 121380 22620 121400
rect 22880 121380 23120 121400
rect 23380 121380 23620 121400
rect 23880 121380 24120 121400
rect 24380 121380 24620 121400
rect 24880 121380 25120 121400
rect 25380 121380 25620 121400
rect 25880 121380 26120 121400
rect 26380 121380 26620 121400
rect 26880 121380 27120 121400
rect 27380 121380 27620 121400
rect 27880 121380 28120 121400
rect 28380 121380 28620 121400
rect 28880 121380 29120 121400
rect 29380 121380 29620 121400
rect 29880 121380 30120 121400
rect 30380 121380 30620 121400
rect 30880 121380 31120 121400
rect 31380 121380 31620 121400
rect 31880 121380 32120 121400
rect 32380 121380 32620 121400
rect 32880 121380 33120 121400
rect 33380 121380 33620 121400
rect 33880 121380 34120 121400
rect 34380 121380 34620 121400
rect 34880 121380 35120 121400
rect 35380 121380 35620 121400
rect 35880 121380 36120 121400
rect 36380 121380 36620 121400
rect 36880 121380 37120 121400
rect 37380 121380 37620 121400
rect 37880 121380 38120 121400
rect 38380 121380 38620 121400
rect 38880 121380 39120 121400
rect 39380 121380 39620 121400
rect 39880 121380 40120 121400
rect 40380 121380 40620 121400
rect 40880 121380 41120 121400
rect 41380 121380 41620 121400
rect 41880 121380 42120 121400
rect 42380 121380 42620 121400
rect 42880 121380 43120 121400
rect 43380 121380 43620 121400
rect 43880 121380 44120 121400
rect 44380 121380 44620 121400
rect 44880 121380 45120 121400
rect 45380 121380 45620 121400
rect 45880 121380 46120 121400
rect 46380 121380 46620 121400
rect 46880 121380 47120 121400
rect 47380 121380 47620 121400
rect 47880 121380 48120 121400
rect 48380 121380 48620 121400
rect 48880 121380 49120 121400
rect 49380 121380 49620 121400
rect 49880 121380 50120 121400
rect 50380 121380 50620 121400
rect 50880 121380 51120 121400
rect 51380 121380 51620 121400
rect 51880 121380 52120 121400
rect 52380 121380 52620 121400
rect 52880 121380 53120 121400
rect 53380 121380 53620 121400
rect 53880 121380 54120 121400
rect 54380 121380 54620 121400
rect 54880 121380 55120 121400
rect 55380 121380 55620 121400
rect 55880 121380 56120 121400
rect 56380 121380 56620 121400
rect 56880 121380 57120 121400
rect 57380 121380 57620 121400
rect 57880 121380 58000 121400
rect 14000 121120 14100 121380
rect 14400 121120 14600 121380
rect 14900 121120 15100 121380
rect 15400 121120 15600 121380
rect 15900 121120 16100 121380
rect 16400 121120 16600 121380
rect 16900 121120 17100 121380
rect 17400 121120 17600 121380
rect 17900 121120 18100 121380
rect 18400 121120 18600 121380
rect 18900 121120 19100 121380
rect 19400 121120 19600 121380
rect 19900 121120 20100 121380
rect 20400 121120 20600 121380
rect 20900 121120 21100 121380
rect 21400 121120 21600 121380
rect 21900 121120 22100 121380
rect 22400 121120 22600 121380
rect 22900 121120 23100 121380
rect 23400 121120 23600 121380
rect 23900 121120 24100 121380
rect 24400 121120 24600 121380
rect 24900 121120 25100 121380
rect 25400 121120 25600 121380
rect 25900 121120 26100 121380
rect 26400 121120 26600 121380
rect 26900 121120 27100 121380
rect 27400 121120 27600 121380
rect 27900 121120 28100 121380
rect 28400 121120 28600 121380
rect 28900 121120 29100 121380
rect 29400 121120 29600 121380
rect 29900 121120 30100 121380
rect 30400 121120 30600 121380
rect 30900 121120 31100 121380
rect 31400 121120 31600 121380
rect 31900 121120 32100 121380
rect 32400 121120 32600 121380
rect 32900 121120 33100 121380
rect 33400 121120 33600 121380
rect 33900 121120 34100 121380
rect 34400 121120 34600 121380
rect 34900 121120 35100 121380
rect 35400 121120 35600 121380
rect 35900 121120 36100 121380
rect 36400 121120 36600 121380
rect 36900 121120 37100 121380
rect 37400 121120 37600 121380
rect 37900 121120 38100 121380
rect 38400 121120 38600 121380
rect 38900 121120 39100 121380
rect 39400 121120 39600 121380
rect 39900 121120 40100 121380
rect 40400 121120 40600 121380
rect 40900 121120 41100 121380
rect 41400 121120 41600 121380
rect 41900 121120 42100 121380
rect 42400 121120 42600 121380
rect 42900 121120 43100 121380
rect 43400 121120 43600 121380
rect 43900 121120 44100 121380
rect 44400 121120 44600 121380
rect 44900 121120 45100 121380
rect 45400 121120 45600 121380
rect 45900 121120 46100 121380
rect 46400 121120 46600 121380
rect 46900 121120 47100 121380
rect 47400 121120 47600 121380
rect 47900 121120 48100 121380
rect 48400 121120 48600 121380
rect 48900 121120 49100 121380
rect 49400 121120 49600 121380
rect 49900 121120 50100 121380
rect 50400 121120 50600 121380
rect 50900 121120 51100 121380
rect 51400 121120 51600 121380
rect 51900 121120 52100 121380
rect 52400 121120 52600 121380
rect 52900 121120 53100 121380
rect 53400 121120 53600 121380
rect 53900 121120 54100 121380
rect 54400 121120 54600 121380
rect 54900 121120 55100 121380
rect 55400 121120 55600 121380
rect 55900 121120 56100 121380
rect 56400 121120 56600 121380
rect 56900 121120 57100 121380
rect 57400 121120 57600 121380
rect 57900 121120 58000 121380
rect 14000 121100 14120 121120
rect 14380 121100 14620 121120
rect 14880 121100 15120 121120
rect 15380 121100 15620 121120
rect 15880 121100 16120 121120
rect 16380 121100 16620 121120
rect 16880 121100 17120 121120
rect 17380 121100 17620 121120
rect 17880 121100 18120 121120
rect 18380 121100 18620 121120
rect 18880 121100 19120 121120
rect 19380 121100 19620 121120
rect 19880 121100 20120 121120
rect 20380 121100 20620 121120
rect 20880 121100 21120 121120
rect 21380 121100 21620 121120
rect 21880 121100 22120 121120
rect 22380 121100 22620 121120
rect 22880 121100 23120 121120
rect 23380 121100 23620 121120
rect 23880 121100 24120 121120
rect 24380 121100 24620 121120
rect 24880 121100 25120 121120
rect 25380 121100 25620 121120
rect 25880 121100 26120 121120
rect 26380 121100 26620 121120
rect 26880 121100 27120 121120
rect 27380 121100 27620 121120
rect 27880 121100 28120 121120
rect 28380 121100 28620 121120
rect 28880 121100 29120 121120
rect 29380 121100 29620 121120
rect 29880 121100 30120 121120
rect 30380 121100 30620 121120
rect 30880 121100 31120 121120
rect 31380 121100 31620 121120
rect 31880 121100 32120 121120
rect 32380 121100 32620 121120
rect 32880 121100 33120 121120
rect 33380 121100 33620 121120
rect 33880 121100 34120 121120
rect 34380 121100 34620 121120
rect 34880 121100 35120 121120
rect 35380 121100 35620 121120
rect 35880 121100 36120 121120
rect 36380 121100 36620 121120
rect 36880 121100 37120 121120
rect 37380 121100 37620 121120
rect 37880 121100 38120 121120
rect 38380 121100 38620 121120
rect 38880 121100 39120 121120
rect 39380 121100 39620 121120
rect 39880 121100 40120 121120
rect 40380 121100 40620 121120
rect 40880 121100 41120 121120
rect 41380 121100 41620 121120
rect 41880 121100 42120 121120
rect 42380 121100 42620 121120
rect 42880 121100 43120 121120
rect 43380 121100 43620 121120
rect 43880 121100 44120 121120
rect 44380 121100 44620 121120
rect 44880 121100 45120 121120
rect 45380 121100 45620 121120
rect 45880 121100 46120 121120
rect 46380 121100 46620 121120
rect 46880 121100 47120 121120
rect 47380 121100 47620 121120
rect 47880 121100 48120 121120
rect 48380 121100 48620 121120
rect 48880 121100 49120 121120
rect 49380 121100 49620 121120
rect 49880 121100 50120 121120
rect 50380 121100 50620 121120
rect 50880 121100 51120 121120
rect 51380 121100 51620 121120
rect 51880 121100 52120 121120
rect 52380 121100 52620 121120
rect 52880 121100 53120 121120
rect 53380 121100 53620 121120
rect 53880 121100 54120 121120
rect 54380 121100 54620 121120
rect 54880 121100 55120 121120
rect 55380 121100 55620 121120
rect 55880 121100 56120 121120
rect 56380 121100 56620 121120
rect 56880 121100 57120 121120
rect 57380 121100 57620 121120
rect 57880 121100 58000 121120
rect 14000 120900 58000 121100
rect 14000 120880 14120 120900
rect 14380 120880 14620 120900
rect 14880 120880 15120 120900
rect 15380 120880 15620 120900
rect 15880 120880 16120 120900
rect 16380 120880 16620 120900
rect 16880 120880 17120 120900
rect 17380 120880 17620 120900
rect 17880 120880 18120 120900
rect 18380 120880 18620 120900
rect 18880 120880 19120 120900
rect 19380 120880 19620 120900
rect 19880 120880 20120 120900
rect 20380 120880 20620 120900
rect 20880 120880 21120 120900
rect 21380 120880 21620 120900
rect 21880 120880 22120 120900
rect 22380 120880 22620 120900
rect 22880 120880 23120 120900
rect 23380 120880 23620 120900
rect 23880 120880 24120 120900
rect 24380 120880 24620 120900
rect 24880 120880 25120 120900
rect 25380 120880 25620 120900
rect 25880 120880 26120 120900
rect 26380 120880 26620 120900
rect 26880 120880 27120 120900
rect 27380 120880 27620 120900
rect 27880 120880 28120 120900
rect 28380 120880 28620 120900
rect 28880 120880 29120 120900
rect 29380 120880 29620 120900
rect 29880 120880 30120 120900
rect 30380 120880 30620 120900
rect 30880 120880 31120 120900
rect 31380 120880 31620 120900
rect 31880 120880 32120 120900
rect 32380 120880 32620 120900
rect 32880 120880 33120 120900
rect 33380 120880 33620 120900
rect 33880 120880 34120 120900
rect 34380 120880 34620 120900
rect 34880 120880 35120 120900
rect 35380 120880 35620 120900
rect 35880 120880 36120 120900
rect 36380 120880 36620 120900
rect 36880 120880 37120 120900
rect 37380 120880 37620 120900
rect 37880 120880 38120 120900
rect 38380 120880 38620 120900
rect 38880 120880 39120 120900
rect 39380 120880 39620 120900
rect 39880 120880 40120 120900
rect 40380 120880 40620 120900
rect 40880 120880 41120 120900
rect 41380 120880 41620 120900
rect 41880 120880 42120 120900
rect 42380 120880 42620 120900
rect 42880 120880 43120 120900
rect 43380 120880 43620 120900
rect 43880 120880 44120 120900
rect 44380 120880 44620 120900
rect 44880 120880 45120 120900
rect 45380 120880 45620 120900
rect 45880 120880 46120 120900
rect 46380 120880 46620 120900
rect 46880 120880 47120 120900
rect 47380 120880 47620 120900
rect 47880 120880 48120 120900
rect 48380 120880 48620 120900
rect 48880 120880 49120 120900
rect 49380 120880 49620 120900
rect 49880 120880 50120 120900
rect 50380 120880 50620 120900
rect 50880 120880 51120 120900
rect 51380 120880 51620 120900
rect 51880 120880 52120 120900
rect 52380 120880 52620 120900
rect 52880 120880 53120 120900
rect 53380 120880 53620 120900
rect 53880 120880 54120 120900
rect 54380 120880 54620 120900
rect 54880 120880 55120 120900
rect 55380 120880 55620 120900
rect 55880 120880 56120 120900
rect 56380 120880 56620 120900
rect 56880 120880 57120 120900
rect 57380 120880 57620 120900
rect 57880 120880 58000 120900
rect 14000 120620 14100 120880
rect 14400 120620 14600 120880
rect 14900 120620 15100 120880
rect 15400 120620 15600 120880
rect 15900 120620 16100 120880
rect 16400 120620 16600 120880
rect 16900 120620 17100 120880
rect 17400 120620 17600 120880
rect 17900 120620 18100 120880
rect 18400 120620 18600 120880
rect 18900 120620 19100 120880
rect 19400 120620 19600 120880
rect 19900 120620 20100 120880
rect 20400 120620 20600 120880
rect 20900 120620 21100 120880
rect 21400 120620 21600 120880
rect 21900 120620 22100 120880
rect 22400 120620 22600 120880
rect 22900 120620 23100 120880
rect 23400 120620 23600 120880
rect 23900 120620 24100 120880
rect 24400 120620 24600 120880
rect 24900 120620 25100 120880
rect 25400 120620 25600 120880
rect 25900 120620 26100 120880
rect 26400 120620 26600 120880
rect 26900 120620 27100 120880
rect 27400 120620 27600 120880
rect 27900 120620 28100 120880
rect 28400 120620 28600 120880
rect 28900 120620 29100 120880
rect 29400 120620 29600 120880
rect 29900 120620 30100 120880
rect 30400 120620 30600 120880
rect 30900 120620 31100 120880
rect 31400 120620 31600 120880
rect 31900 120620 32100 120880
rect 32400 120620 32600 120880
rect 32900 120620 33100 120880
rect 33400 120620 33600 120880
rect 33900 120620 34100 120880
rect 34400 120620 34600 120880
rect 34900 120620 35100 120880
rect 35400 120620 35600 120880
rect 35900 120620 36100 120880
rect 36400 120620 36600 120880
rect 36900 120620 37100 120880
rect 37400 120620 37600 120880
rect 37900 120620 38100 120880
rect 38400 120620 38600 120880
rect 38900 120620 39100 120880
rect 39400 120620 39600 120880
rect 39900 120620 40100 120880
rect 40400 120620 40600 120880
rect 40900 120620 41100 120880
rect 41400 120620 41600 120880
rect 41900 120620 42100 120880
rect 42400 120620 42600 120880
rect 42900 120620 43100 120880
rect 43400 120620 43600 120880
rect 43900 120620 44100 120880
rect 44400 120620 44600 120880
rect 44900 120620 45100 120880
rect 45400 120620 45600 120880
rect 45900 120620 46100 120880
rect 46400 120620 46600 120880
rect 46900 120620 47100 120880
rect 47400 120620 47600 120880
rect 47900 120620 48100 120880
rect 48400 120620 48600 120880
rect 48900 120620 49100 120880
rect 49400 120620 49600 120880
rect 49900 120620 50100 120880
rect 50400 120620 50600 120880
rect 50900 120620 51100 120880
rect 51400 120620 51600 120880
rect 51900 120620 52100 120880
rect 52400 120620 52600 120880
rect 52900 120620 53100 120880
rect 53400 120620 53600 120880
rect 53900 120620 54100 120880
rect 54400 120620 54600 120880
rect 54900 120620 55100 120880
rect 55400 120620 55600 120880
rect 55900 120620 56100 120880
rect 56400 120620 56600 120880
rect 56900 120620 57100 120880
rect 57400 120620 57600 120880
rect 57900 120620 58000 120880
rect 14000 120600 14120 120620
rect 14380 120600 14620 120620
rect 14880 120600 15120 120620
rect 15380 120600 15620 120620
rect 15880 120600 16120 120620
rect 16380 120600 16620 120620
rect 16880 120600 17120 120620
rect 17380 120600 17620 120620
rect 17880 120600 18120 120620
rect 18380 120600 18620 120620
rect 18880 120600 19120 120620
rect 19380 120600 19620 120620
rect 19880 120600 20120 120620
rect 20380 120600 20620 120620
rect 20880 120600 21120 120620
rect 21380 120600 21620 120620
rect 21880 120600 22120 120620
rect 22380 120600 22620 120620
rect 22880 120600 23120 120620
rect 23380 120600 23620 120620
rect 23880 120600 24120 120620
rect 24380 120600 24620 120620
rect 24880 120600 25120 120620
rect 25380 120600 25620 120620
rect 25880 120600 26120 120620
rect 26380 120600 26620 120620
rect 26880 120600 27120 120620
rect 27380 120600 27620 120620
rect 27880 120600 28120 120620
rect 28380 120600 28620 120620
rect 28880 120600 29120 120620
rect 29380 120600 29620 120620
rect 29880 120600 30120 120620
rect 30380 120600 30620 120620
rect 30880 120600 31120 120620
rect 31380 120600 31620 120620
rect 31880 120600 32120 120620
rect 32380 120600 32620 120620
rect 32880 120600 33120 120620
rect 33380 120600 33620 120620
rect 33880 120600 34120 120620
rect 34380 120600 34620 120620
rect 34880 120600 35120 120620
rect 35380 120600 35620 120620
rect 35880 120600 36120 120620
rect 36380 120600 36620 120620
rect 36880 120600 37120 120620
rect 37380 120600 37620 120620
rect 37880 120600 38120 120620
rect 38380 120600 38620 120620
rect 38880 120600 39120 120620
rect 39380 120600 39620 120620
rect 39880 120600 40120 120620
rect 40380 120600 40620 120620
rect 40880 120600 41120 120620
rect 41380 120600 41620 120620
rect 41880 120600 42120 120620
rect 42380 120600 42620 120620
rect 42880 120600 43120 120620
rect 43380 120600 43620 120620
rect 43880 120600 44120 120620
rect 44380 120600 44620 120620
rect 44880 120600 45120 120620
rect 45380 120600 45620 120620
rect 45880 120600 46120 120620
rect 46380 120600 46620 120620
rect 46880 120600 47120 120620
rect 47380 120600 47620 120620
rect 47880 120600 48120 120620
rect 48380 120600 48620 120620
rect 48880 120600 49120 120620
rect 49380 120600 49620 120620
rect 49880 120600 50120 120620
rect 50380 120600 50620 120620
rect 50880 120600 51120 120620
rect 51380 120600 51620 120620
rect 51880 120600 52120 120620
rect 52380 120600 52620 120620
rect 52880 120600 53120 120620
rect 53380 120600 53620 120620
rect 53880 120600 54120 120620
rect 54380 120600 54620 120620
rect 54880 120600 55120 120620
rect 55380 120600 55620 120620
rect 55880 120600 56120 120620
rect 56380 120600 56620 120620
rect 56880 120600 57120 120620
rect 57380 120600 57620 120620
rect 57880 120600 58000 120620
rect 14000 120400 58000 120600
rect 14000 120380 14120 120400
rect 14380 120380 14620 120400
rect 14880 120380 15120 120400
rect 15380 120380 15620 120400
rect 15880 120380 16120 120400
rect 16380 120380 16620 120400
rect 16880 120380 17120 120400
rect 17380 120380 17620 120400
rect 17880 120380 18120 120400
rect 18380 120380 18620 120400
rect 18880 120380 19120 120400
rect 19380 120380 19620 120400
rect 19880 120380 20120 120400
rect 20380 120380 20620 120400
rect 20880 120380 21120 120400
rect 21380 120380 21620 120400
rect 21880 120380 22120 120400
rect 22380 120380 22620 120400
rect 22880 120380 23120 120400
rect 23380 120380 23620 120400
rect 23880 120380 24120 120400
rect 24380 120380 24620 120400
rect 24880 120380 25120 120400
rect 25380 120380 25620 120400
rect 25880 120380 26120 120400
rect 26380 120380 26620 120400
rect 26880 120380 27120 120400
rect 27380 120380 27620 120400
rect 27880 120380 28120 120400
rect 28380 120380 28620 120400
rect 28880 120380 29120 120400
rect 29380 120380 29620 120400
rect 29880 120380 30120 120400
rect 30380 120380 30620 120400
rect 30880 120380 31120 120400
rect 31380 120380 31620 120400
rect 31880 120380 32120 120400
rect 32380 120380 32620 120400
rect 32880 120380 33120 120400
rect 33380 120380 33620 120400
rect 33880 120380 34120 120400
rect 34380 120380 34620 120400
rect 34880 120380 35120 120400
rect 35380 120380 35620 120400
rect 35880 120380 36120 120400
rect 36380 120380 36620 120400
rect 36880 120380 37120 120400
rect 37380 120380 37620 120400
rect 37880 120380 38120 120400
rect 38380 120380 38620 120400
rect 38880 120380 39120 120400
rect 39380 120380 39620 120400
rect 39880 120380 40120 120400
rect 40380 120380 40620 120400
rect 40880 120380 41120 120400
rect 41380 120380 41620 120400
rect 41880 120380 42120 120400
rect 42380 120380 42620 120400
rect 42880 120380 43120 120400
rect 43380 120380 43620 120400
rect 43880 120380 44120 120400
rect 44380 120380 44620 120400
rect 44880 120380 45120 120400
rect 45380 120380 45620 120400
rect 45880 120380 46120 120400
rect 46380 120380 46620 120400
rect 46880 120380 47120 120400
rect 47380 120380 47620 120400
rect 47880 120380 48120 120400
rect 48380 120380 48620 120400
rect 48880 120380 49120 120400
rect 49380 120380 49620 120400
rect 49880 120380 50120 120400
rect 50380 120380 50620 120400
rect 50880 120380 51120 120400
rect 51380 120380 51620 120400
rect 51880 120380 52120 120400
rect 52380 120380 52620 120400
rect 52880 120380 53120 120400
rect 53380 120380 53620 120400
rect 53880 120380 54120 120400
rect 54380 120380 54620 120400
rect 54880 120380 55120 120400
rect 55380 120380 55620 120400
rect 55880 120380 56120 120400
rect 56380 120380 56620 120400
rect 56880 120380 57120 120400
rect 57380 120380 57620 120400
rect 57880 120380 58000 120400
rect 14000 120120 14100 120380
rect 14400 120120 14600 120380
rect 14900 120120 15100 120380
rect 15400 120120 15600 120380
rect 15900 120120 16100 120380
rect 16400 120120 16600 120380
rect 16900 120120 17100 120380
rect 17400 120120 17600 120380
rect 17900 120120 18100 120380
rect 18400 120120 18600 120380
rect 18900 120120 19100 120380
rect 19400 120120 19600 120380
rect 19900 120120 20100 120380
rect 20400 120120 20600 120380
rect 20900 120120 21100 120380
rect 21400 120120 21600 120380
rect 21900 120120 22100 120380
rect 22400 120120 22600 120380
rect 22900 120120 23100 120380
rect 23400 120120 23600 120380
rect 23900 120120 24100 120380
rect 24400 120120 24600 120380
rect 24900 120120 25100 120380
rect 25400 120120 25600 120380
rect 25900 120120 26100 120380
rect 26400 120120 26600 120380
rect 26900 120120 27100 120380
rect 27400 120120 27600 120380
rect 27900 120120 28100 120380
rect 28400 120120 28600 120380
rect 28900 120120 29100 120380
rect 29400 120120 29600 120380
rect 29900 120120 30100 120380
rect 30400 120120 30600 120380
rect 30900 120120 31100 120380
rect 31400 120120 31600 120380
rect 31900 120120 32100 120380
rect 32400 120120 32600 120380
rect 32900 120120 33100 120380
rect 33400 120120 33600 120380
rect 33900 120120 34100 120380
rect 34400 120120 34600 120380
rect 34900 120120 35100 120380
rect 35400 120120 35600 120380
rect 35900 120120 36100 120380
rect 36400 120120 36600 120380
rect 36900 120120 37100 120380
rect 37400 120120 37600 120380
rect 37900 120120 38100 120380
rect 38400 120120 38600 120380
rect 38900 120120 39100 120380
rect 39400 120120 39600 120380
rect 39900 120120 40100 120380
rect 40400 120120 40600 120380
rect 40900 120120 41100 120380
rect 41400 120120 41600 120380
rect 41900 120120 42100 120380
rect 42400 120120 42600 120380
rect 42900 120120 43100 120380
rect 43400 120120 43600 120380
rect 43900 120120 44100 120380
rect 44400 120120 44600 120380
rect 44900 120120 45100 120380
rect 45400 120120 45600 120380
rect 45900 120120 46100 120380
rect 46400 120120 46600 120380
rect 46900 120120 47100 120380
rect 47400 120120 47600 120380
rect 47900 120120 48100 120380
rect 48400 120120 48600 120380
rect 48900 120120 49100 120380
rect 49400 120120 49600 120380
rect 49900 120120 50100 120380
rect 50400 120120 50600 120380
rect 50900 120120 51100 120380
rect 51400 120120 51600 120380
rect 51900 120120 52100 120380
rect 52400 120120 52600 120380
rect 52900 120120 53100 120380
rect 53400 120120 53600 120380
rect 53900 120120 54100 120380
rect 54400 120120 54600 120380
rect 54900 120120 55100 120380
rect 55400 120120 55600 120380
rect 55900 120120 56100 120380
rect 56400 120120 56600 120380
rect 56900 120120 57100 120380
rect 57400 120120 57600 120380
rect 57900 120120 58000 120380
rect 14000 120100 14120 120120
rect 14380 120100 14620 120120
rect 14880 120100 15120 120120
rect 15380 120100 15620 120120
rect 15880 120100 16120 120120
rect 16380 120100 16620 120120
rect 16880 120100 17120 120120
rect 17380 120100 17620 120120
rect 17880 120100 18120 120120
rect 18380 120100 18620 120120
rect 18880 120100 19120 120120
rect 19380 120100 19620 120120
rect 19880 120100 20120 120120
rect 20380 120100 20620 120120
rect 20880 120100 21120 120120
rect 21380 120100 21620 120120
rect 21880 120100 22120 120120
rect 22380 120100 22620 120120
rect 22880 120100 23120 120120
rect 23380 120100 23620 120120
rect 23880 120100 24120 120120
rect 24380 120100 24620 120120
rect 24880 120100 25120 120120
rect 25380 120100 25620 120120
rect 25880 120100 26120 120120
rect 26380 120100 26620 120120
rect 26880 120100 27120 120120
rect 27380 120100 27620 120120
rect 27880 120100 28120 120120
rect 28380 120100 28620 120120
rect 28880 120100 29120 120120
rect 29380 120100 29620 120120
rect 29880 120100 30120 120120
rect 30380 120100 30620 120120
rect 30880 120100 31120 120120
rect 31380 120100 31620 120120
rect 31880 120100 32120 120120
rect 32380 120100 32620 120120
rect 32880 120100 33120 120120
rect 33380 120100 33620 120120
rect 33880 120100 34120 120120
rect 34380 120100 34620 120120
rect 34880 120100 35120 120120
rect 35380 120100 35620 120120
rect 35880 120100 36120 120120
rect 36380 120100 36620 120120
rect 36880 120100 37120 120120
rect 37380 120100 37620 120120
rect 37880 120100 38120 120120
rect 38380 120100 38620 120120
rect 38880 120100 39120 120120
rect 39380 120100 39620 120120
rect 39880 120100 40120 120120
rect 40380 120100 40620 120120
rect 40880 120100 41120 120120
rect 41380 120100 41620 120120
rect 41880 120100 42120 120120
rect 42380 120100 42620 120120
rect 42880 120100 43120 120120
rect 43380 120100 43620 120120
rect 43880 120100 44120 120120
rect 44380 120100 44620 120120
rect 44880 120100 45120 120120
rect 45380 120100 45620 120120
rect 45880 120100 46120 120120
rect 46380 120100 46620 120120
rect 46880 120100 47120 120120
rect 47380 120100 47620 120120
rect 47880 120100 48120 120120
rect 48380 120100 48620 120120
rect 48880 120100 49120 120120
rect 49380 120100 49620 120120
rect 49880 120100 50120 120120
rect 50380 120100 50620 120120
rect 50880 120100 51120 120120
rect 51380 120100 51620 120120
rect 51880 120100 52120 120120
rect 52380 120100 52620 120120
rect 52880 120100 53120 120120
rect 53380 120100 53620 120120
rect 53880 120100 54120 120120
rect 54380 120100 54620 120120
rect 54880 120100 55120 120120
rect 55380 120100 55620 120120
rect 55880 120100 56120 120120
rect 56380 120100 56620 120120
rect 56880 120100 57120 120120
rect 57380 120100 57620 120120
rect 57880 120100 58000 120120
rect 14000 119900 58000 120100
rect 14000 119880 14120 119900
rect 14380 119880 14620 119900
rect 14880 119880 15120 119900
rect 15380 119880 15620 119900
rect 15880 119880 16120 119900
rect 16380 119880 16620 119900
rect 16880 119880 17120 119900
rect 17380 119880 17620 119900
rect 17880 119880 18120 119900
rect 18380 119880 18620 119900
rect 18880 119880 19120 119900
rect 19380 119880 19620 119900
rect 19880 119880 20120 119900
rect 20380 119880 20620 119900
rect 20880 119880 21120 119900
rect 21380 119880 21620 119900
rect 21880 119880 22120 119900
rect 22380 119880 22620 119900
rect 22880 119880 23120 119900
rect 23380 119880 23620 119900
rect 23880 119880 24120 119900
rect 24380 119880 24620 119900
rect 24880 119880 25120 119900
rect 25380 119880 25620 119900
rect 25880 119880 26120 119900
rect 26380 119880 26620 119900
rect 26880 119880 27120 119900
rect 27380 119880 27620 119900
rect 27880 119880 28120 119900
rect 28380 119880 28620 119900
rect 28880 119880 29120 119900
rect 29380 119880 29620 119900
rect 29880 119880 30120 119900
rect 30380 119880 30620 119900
rect 30880 119880 31120 119900
rect 31380 119880 31620 119900
rect 31880 119880 32120 119900
rect 32380 119880 32620 119900
rect 32880 119880 33120 119900
rect 33380 119880 33620 119900
rect 33880 119880 34120 119900
rect 34380 119880 34620 119900
rect 34880 119880 35120 119900
rect 35380 119880 35620 119900
rect 35880 119880 36120 119900
rect 36380 119880 36620 119900
rect 36880 119880 37120 119900
rect 37380 119880 37620 119900
rect 37880 119880 38120 119900
rect 38380 119880 38620 119900
rect 38880 119880 39120 119900
rect 39380 119880 39620 119900
rect 39880 119880 40120 119900
rect 40380 119880 40620 119900
rect 40880 119880 41120 119900
rect 41380 119880 41620 119900
rect 41880 119880 42120 119900
rect 42380 119880 42620 119900
rect 42880 119880 43120 119900
rect 43380 119880 43620 119900
rect 43880 119880 44120 119900
rect 44380 119880 44620 119900
rect 44880 119880 45120 119900
rect 45380 119880 45620 119900
rect 45880 119880 46120 119900
rect 46380 119880 46620 119900
rect 46880 119880 47120 119900
rect 47380 119880 47620 119900
rect 47880 119880 48120 119900
rect 48380 119880 48620 119900
rect 48880 119880 49120 119900
rect 49380 119880 49620 119900
rect 49880 119880 50120 119900
rect 50380 119880 50620 119900
rect 50880 119880 51120 119900
rect 51380 119880 51620 119900
rect 51880 119880 52120 119900
rect 52380 119880 52620 119900
rect 52880 119880 53120 119900
rect 53380 119880 53620 119900
rect 53880 119880 54120 119900
rect 54380 119880 54620 119900
rect 54880 119880 55120 119900
rect 55380 119880 55620 119900
rect 55880 119880 56120 119900
rect 56380 119880 56620 119900
rect 56880 119880 57120 119900
rect 57380 119880 57620 119900
rect 57880 119880 58000 119900
rect 14000 119620 14100 119880
rect 14400 119620 14600 119880
rect 14900 119620 15100 119880
rect 15400 119620 15600 119880
rect 15900 119620 16100 119880
rect 16400 119620 16600 119880
rect 16900 119620 17100 119880
rect 17400 119620 17600 119880
rect 17900 119620 18100 119880
rect 18400 119620 18600 119880
rect 18900 119620 19100 119880
rect 19400 119620 19600 119880
rect 19900 119620 20100 119880
rect 20400 119620 20600 119880
rect 20900 119620 21100 119880
rect 21400 119620 21600 119880
rect 21900 119620 22100 119880
rect 22400 119620 22600 119880
rect 22900 119620 23100 119880
rect 23400 119620 23600 119880
rect 23900 119620 24100 119880
rect 24400 119620 24600 119880
rect 24900 119620 25100 119880
rect 25400 119620 25600 119880
rect 25900 119620 26100 119880
rect 26400 119620 26600 119880
rect 26900 119620 27100 119880
rect 27400 119620 27600 119880
rect 27900 119620 28100 119880
rect 28400 119620 28600 119880
rect 28900 119620 29100 119880
rect 29400 119620 29600 119880
rect 29900 119620 30100 119880
rect 30400 119620 30600 119880
rect 30900 119620 31100 119880
rect 31400 119620 31600 119880
rect 31900 119620 32100 119880
rect 32400 119620 32600 119880
rect 32900 119620 33100 119880
rect 33400 119620 33600 119880
rect 33900 119620 34100 119880
rect 34400 119620 34600 119880
rect 34900 119620 35100 119880
rect 35400 119620 35600 119880
rect 35900 119620 36100 119880
rect 36400 119620 36600 119880
rect 36900 119620 37100 119880
rect 37400 119620 37600 119880
rect 37900 119620 38100 119880
rect 38400 119620 38600 119880
rect 38900 119620 39100 119880
rect 39400 119620 39600 119880
rect 39900 119620 40100 119880
rect 40400 119620 40600 119880
rect 40900 119620 41100 119880
rect 41400 119620 41600 119880
rect 41900 119620 42100 119880
rect 42400 119620 42600 119880
rect 42900 119620 43100 119880
rect 43400 119620 43600 119880
rect 43900 119620 44100 119880
rect 44400 119620 44600 119880
rect 44900 119620 45100 119880
rect 45400 119620 45600 119880
rect 45900 119620 46100 119880
rect 46400 119620 46600 119880
rect 46900 119620 47100 119880
rect 47400 119620 47600 119880
rect 47900 119620 48100 119880
rect 48400 119620 48600 119880
rect 48900 119620 49100 119880
rect 49400 119620 49600 119880
rect 49900 119620 50100 119880
rect 50400 119620 50600 119880
rect 50900 119620 51100 119880
rect 51400 119620 51600 119880
rect 51900 119620 52100 119880
rect 52400 119620 52600 119880
rect 52900 119620 53100 119880
rect 53400 119620 53600 119880
rect 53900 119620 54100 119880
rect 54400 119620 54600 119880
rect 54900 119620 55100 119880
rect 55400 119620 55600 119880
rect 55900 119620 56100 119880
rect 56400 119620 56600 119880
rect 56900 119620 57100 119880
rect 57400 119620 57600 119880
rect 57900 119620 58000 119880
rect 14000 119600 14120 119620
rect 14380 119600 14620 119620
rect 14880 119600 15120 119620
rect 15380 119600 15620 119620
rect 15880 119600 16120 119620
rect 16380 119600 16620 119620
rect 16880 119600 17120 119620
rect 17380 119600 17620 119620
rect 17880 119600 18120 119620
rect 18380 119600 18620 119620
rect 18880 119600 19120 119620
rect 19380 119600 19620 119620
rect 19880 119600 20120 119620
rect 20380 119600 20620 119620
rect 20880 119600 21120 119620
rect 21380 119600 21620 119620
rect 21880 119600 22120 119620
rect 22380 119600 22620 119620
rect 22880 119600 23120 119620
rect 23380 119600 23620 119620
rect 23880 119600 24120 119620
rect 24380 119600 24620 119620
rect 24880 119600 25120 119620
rect 25380 119600 25620 119620
rect 25880 119600 26120 119620
rect 26380 119600 26620 119620
rect 26880 119600 27120 119620
rect 27380 119600 27620 119620
rect 27880 119600 28120 119620
rect 28380 119600 28620 119620
rect 28880 119600 29120 119620
rect 29380 119600 29620 119620
rect 29880 119600 30120 119620
rect 30380 119600 30620 119620
rect 30880 119600 31120 119620
rect 31380 119600 31620 119620
rect 31880 119600 32120 119620
rect 32380 119600 32620 119620
rect 32880 119600 33120 119620
rect 33380 119600 33620 119620
rect 33880 119600 34120 119620
rect 34380 119600 34620 119620
rect 34880 119600 35120 119620
rect 35380 119600 35620 119620
rect 35880 119600 36120 119620
rect 36380 119600 36620 119620
rect 36880 119600 37120 119620
rect 37380 119600 37620 119620
rect 37880 119600 38120 119620
rect 38380 119600 38620 119620
rect 38880 119600 39120 119620
rect 39380 119600 39620 119620
rect 39880 119600 40120 119620
rect 40380 119600 40620 119620
rect 40880 119600 41120 119620
rect 41380 119600 41620 119620
rect 41880 119600 42120 119620
rect 42380 119600 42620 119620
rect 42880 119600 43120 119620
rect 43380 119600 43620 119620
rect 43880 119600 44120 119620
rect 44380 119600 44620 119620
rect 44880 119600 45120 119620
rect 45380 119600 45620 119620
rect 45880 119600 46120 119620
rect 46380 119600 46620 119620
rect 46880 119600 47120 119620
rect 47380 119600 47620 119620
rect 47880 119600 48120 119620
rect 48380 119600 48620 119620
rect 48880 119600 49120 119620
rect 49380 119600 49620 119620
rect 49880 119600 50120 119620
rect 50380 119600 50620 119620
rect 50880 119600 51120 119620
rect 51380 119600 51620 119620
rect 51880 119600 52120 119620
rect 52380 119600 52620 119620
rect 52880 119600 53120 119620
rect 53380 119600 53620 119620
rect 53880 119600 54120 119620
rect 54380 119600 54620 119620
rect 54880 119600 55120 119620
rect 55380 119600 55620 119620
rect 55880 119600 56120 119620
rect 56380 119600 56620 119620
rect 56880 119600 57120 119620
rect 57380 119600 57620 119620
rect 57880 119600 58000 119620
rect 14000 119400 58000 119600
rect 14000 119380 14120 119400
rect 14380 119380 14620 119400
rect 14880 119380 15120 119400
rect 15380 119380 15620 119400
rect 15880 119380 16120 119400
rect 16380 119380 16620 119400
rect 16880 119380 17120 119400
rect 17380 119380 17620 119400
rect 17880 119380 18120 119400
rect 18380 119380 18620 119400
rect 18880 119380 19120 119400
rect 19380 119380 19620 119400
rect 19880 119380 20120 119400
rect 20380 119380 20620 119400
rect 20880 119380 21120 119400
rect 21380 119380 21620 119400
rect 21880 119380 22120 119400
rect 22380 119380 22620 119400
rect 22880 119380 23120 119400
rect 23380 119380 23620 119400
rect 23880 119380 24120 119400
rect 24380 119380 24620 119400
rect 24880 119380 25120 119400
rect 25380 119380 25620 119400
rect 25880 119380 26120 119400
rect 26380 119380 26620 119400
rect 26880 119380 27120 119400
rect 27380 119380 27620 119400
rect 27880 119380 28120 119400
rect 28380 119380 28620 119400
rect 28880 119380 29120 119400
rect 29380 119380 29620 119400
rect 29880 119380 30120 119400
rect 30380 119380 30620 119400
rect 30880 119380 31120 119400
rect 31380 119380 31620 119400
rect 31880 119380 32120 119400
rect 32380 119380 32620 119400
rect 32880 119380 33120 119400
rect 33380 119380 33620 119400
rect 33880 119380 34120 119400
rect 34380 119380 34620 119400
rect 34880 119380 35120 119400
rect 35380 119380 35620 119400
rect 35880 119380 36120 119400
rect 36380 119380 36620 119400
rect 36880 119380 37120 119400
rect 37380 119380 37620 119400
rect 37880 119380 38120 119400
rect 38380 119380 38620 119400
rect 38880 119380 39120 119400
rect 39380 119380 39620 119400
rect 39880 119380 40120 119400
rect 40380 119380 40620 119400
rect 40880 119380 41120 119400
rect 41380 119380 41620 119400
rect 41880 119380 42120 119400
rect 42380 119380 42620 119400
rect 42880 119380 43120 119400
rect 43380 119380 43620 119400
rect 43880 119380 44120 119400
rect 44380 119380 44620 119400
rect 44880 119380 45120 119400
rect 45380 119380 45620 119400
rect 45880 119380 46120 119400
rect 46380 119380 46620 119400
rect 46880 119380 47120 119400
rect 47380 119380 47620 119400
rect 47880 119380 48120 119400
rect 48380 119380 48620 119400
rect 48880 119380 49120 119400
rect 49380 119380 49620 119400
rect 49880 119380 50120 119400
rect 50380 119380 50620 119400
rect 50880 119380 51120 119400
rect 51380 119380 51620 119400
rect 51880 119380 52120 119400
rect 52380 119380 52620 119400
rect 52880 119380 53120 119400
rect 53380 119380 53620 119400
rect 53880 119380 54120 119400
rect 54380 119380 54620 119400
rect 54880 119380 55120 119400
rect 55380 119380 55620 119400
rect 55880 119380 56120 119400
rect 56380 119380 56620 119400
rect 56880 119380 57120 119400
rect 57380 119380 57620 119400
rect 57880 119380 58000 119400
rect 14000 119120 14100 119380
rect 14400 119120 14600 119380
rect 14900 119120 15100 119380
rect 15400 119120 15600 119380
rect 15900 119120 16100 119380
rect 16400 119120 16600 119380
rect 16900 119120 17100 119380
rect 17400 119120 17600 119380
rect 17900 119120 18100 119380
rect 18400 119120 18600 119380
rect 18900 119120 19100 119380
rect 19400 119120 19600 119380
rect 19900 119120 20100 119380
rect 20400 119120 20600 119380
rect 20900 119120 21100 119380
rect 21400 119120 21600 119380
rect 21900 119120 22100 119380
rect 22400 119120 22600 119380
rect 22900 119120 23100 119380
rect 23400 119120 23600 119380
rect 23900 119120 24100 119380
rect 24400 119120 24600 119380
rect 24900 119120 25100 119380
rect 25400 119120 25600 119380
rect 25900 119120 26100 119380
rect 26400 119120 26600 119380
rect 26900 119120 27100 119380
rect 27400 119120 27600 119380
rect 27900 119120 28100 119380
rect 28400 119120 28600 119380
rect 28900 119120 29100 119380
rect 29400 119120 29600 119380
rect 29900 119120 30100 119380
rect 30400 119120 30600 119380
rect 30900 119120 31100 119380
rect 31400 119120 31600 119380
rect 31900 119120 32100 119380
rect 32400 119120 32600 119380
rect 32900 119120 33100 119380
rect 33400 119120 33600 119380
rect 33900 119120 34100 119380
rect 34400 119120 34600 119380
rect 34900 119120 35100 119380
rect 35400 119120 35600 119380
rect 35900 119120 36100 119380
rect 36400 119120 36600 119380
rect 36900 119120 37100 119380
rect 37400 119120 37600 119380
rect 37900 119120 38100 119380
rect 38400 119120 38600 119380
rect 38900 119120 39100 119380
rect 39400 119120 39600 119380
rect 39900 119120 40100 119380
rect 40400 119120 40600 119380
rect 40900 119120 41100 119380
rect 41400 119120 41600 119380
rect 41900 119120 42100 119380
rect 42400 119120 42600 119380
rect 42900 119120 43100 119380
rect 43400 119120 43600 119380
rect 43900 119120 44100 119380
rect 44400 119120 44600 119380
rect 44900 119120 45100 119380
rect 45400 119120 45600 119380
rect 45900 119120 46100 119380
rect 46400 119120 46600 119380
rect 46900 119120 47100 119380
rect 47400 119120 47600 119380
rect 47900 119120 48100 119380
rect 48400 119120 48600 119380
rect 48900 119120 49100 119380
rect 49400 119120 49600 119380
rect 49900 119120 50100 119380
rect 50400 119120 50600 119380
rect 50900 119120 51100 119380
rect 51400 119120 51600 119380
rect 51900 119120 52100 119380
rect 52400 119120 52600 119380
rect 52900 119120 53100 119380
rect 53400 119120 53600 119380
rect 53900 119120 54100 119380
rect 54400 119120 54600 119380
rect 54900 119120 55100 119380
rect 55400 119120 55600 119380
rect 55900 119120 56100 119380
rect 56400 119120 56600 119380
rect 56900 119120 57100 119380
rect 57400 119120 57600 119380
rect 57900 119120 58000 119380
rect 14000 119100 14120 119120
rect 14380 119100 14620 119120
rect 14880 119100 15120 119120
rect 15380 119100 15620 119120
rect 15880 119100 16120 119120
rect 16380 119100 16620 119120
rect 16880 119100 17120 119120
rect 17380 119100 17620 119120
rect 17880 119100 18120 119120
rect 18380 119100 18620 119120
rect 18880 119100 19120 119120
rect 19380 119100 19620 119120
rect 19880 119100 20120 119120
rect 20380 119100 20620 119120
rect 20880 119100 21120 119120
rect 21380 119100 21620 119120
rect 21880 119100 22120 119120
rect 22380 119100 22620 119120
rect 22880 119100 23120 119120
rect 23380 119100 23620 119120
rect 23880 119100 24120 119120
rect 24380 119100 24620 119120
rect 24880 119100 25120 119120
rect 25380 119100 25620 119120
rect 25880 119100 26120 119120
rect 26380 119100 26620 119120
rect 26880 119100 27120 119120
rect 27380 119100 27620 119120
rect 27880 119100 28120 119120
rect 28380 119100 28620 119120
rect 28880 119100 29120 119120
rect 29380 119100 29620 119120
rect 29880 119100 30120 119120
rect 30380 119100 30620 119120
rect 30880 119100 31120 119120
rect 31380 119100 31620 119120
rect 31880 119100 32120 119120
rect 32380 119100 32620 119120
rect 32880 119100 33120 119120
rect 33380 119100 33620 119120
rect 33880 119100 34120 119120
rect 34380 119100 34620 119120
rect 34880 119100 35120 119120
rect 35380 119100 35620 119120
rect 35880 119100 36120 119120
rect 36380 119100 36620 119120
rect 36880 119100 37120 119120
rect 37380 119100 37620 119120
rect 37880 119100 38120 119120
rect 38380 119100 38620 119120
rect 38880 119100 39120 119120
rect 39380 119100 39620 119120
rect 39880 119100 40120 119120
rect 40380 119100 40620 119120
rect 40880 119100 41120 119120
rect 41380 119100 41620 119120
rect 41880 119100 42120 119120
rect 42380 119100 42620 119120
rect 42880 119100 43120 119120
rect 43380 119100 43620 119120
rect 43880 119100 44120 119120
rect 44380 119100 44620 119120
rect 44880 119100 45120 119120
rect 45380 119100 45620 119120
rect 45880 119100 46120 119120
rect 46380 119100 46620 119120
rect 46880 119100 47120 119120
rect 47380 119100 47620 119120
rect 47880 119100 48120 119120
rect 48380 119100 48620 119120
rect 48880 119100 49120 119120
rect 49380 119100 49620 119120
rect 49880 119100 50120 119120
rect 50380 119100 50620 119120
rect 50880 119100 51120 119120
rect 51380 119100 51620 119120
rect 51880 119100 52120 119120
rect 52380 119100 52620 119120
rect 52880 119100 53120 119120
rect 53380 119100 53620 119120
rect 53880 119100 54120 119120
rect 54380 119100 54620 119120
rect 54880 119100 55120 119120
rect 55380 119100 55620 119120
rect 55880 119100 56120 119120
rect 56380 119100 56620 119120
rect 56880 119100 57120 119120
rect 57380 119100 57620 119120
rect 57880 119100 58000 119120
rect 14000 118900 58000 119100
rect 14000 118880 14120 118900
rect 14380 118880 14620 118900
rect 14880 118880 15120 118900
rect 15380 118880 15620 118900
rect 15880 118880 16120 118900
rect 16380 118880 16620 118900
rect 16880 118880 17120 118900
rect 17380 118880 17620 118900
rect 17880 118880 18120 118900
rect 18380 118880 18620 118900
rect 18880 118880 19120 118900
rect 19380 118880 19620 118900
rect 19880 118880 20120 118900
rect 20380 118880 20620 118900
rect 20880 118880 21120 118900
rect 21380 118880 21620 118900
rect 21880 118880 22120 118900
rect 22380 118880 22620 118900
rect 22880 118880 23120 118900
rect 23380 118880 23620 118900
rect 23880 118880 24120 118900
rect 24380 118880 24620 118900
rect 24880 118880 25120 118900
rect 25380 118880 25620 118900
rect 25880 118880 26120 118900
rect 26380 118880 26620 118900
rect 26880 118880 27120 118900
rect 27380 118880 27620 118900
rect 27880 118880 28120 118900
rect 28380 118880 28620 118900
rect 28880 118880 29120 118900
rect 29380 118880 29620 118900
rect 29880 118880 30120 118900
rect 30380 118880 30620 118900
rect 30880 118880 31120 118900
rect 31380 118880 31620 118900
rect 31880 118880 32120 118900
rect 32380 118880 32620 118900
rect 32880 118880 33120 118900
rect 33380 118880 33620 118900
rect 33880 118880 34120 118900
rect 34380 118880 34620 118900
rect 34880 118880 35120 118900
rect 35380 118880 35620 118900
rect 35880 118880 36120 118900
rect 36380 118880 36620 118900
rect 36880 118880 37120 118900
rect 37380 118880 37620 118900
rect 37880 118880 38120 118900
rect 38380 118880 38620 118900
rect 38880 118880 39120 118900
rect 39380 118880 39620 118900
rect 39880 118880 40120 118900
rect 40380 118880 40620 118900
rect 40880 118880 41120 118900
rect 41380 118880 41620 118900
rect 41880 118880 42120 118900
rect 42380 118880 42620 118900
rect 42880 118880 43120 118900
rect 43380 118880 43620 118900
rect 43880 118880 44120 118900
rect 44380 118880 44620 118900
rect 44880 118880 45120 118900
rect 45380 118880 45620 118900
rect 45880 118880 46120 118900
rect 46380 118880 46620 118900
rect 46880 118880 47120 118900
rect 47380 118880 47620 118900
rect 47880 118880 48120 118900
rect 48380 118880 48620 118900
rect 48880 118880 49120 118900
rect 49380 118880 49620 118900
rect 49880 118880 50120 118900
rect 50380 118880 50620 118900
rect 50880 118880 51120 118900
rect 51380 118880 51620 118900
rect 51880 118880 52120 118900
rect 52380 118880 52620 118900
rect 52880 118880 53120 118900
rect 53380 118880 53620 118900
rect 53880 118880 54120 118900
rect 54380 118880 54620 118900
rect 54880 118880 55120 118900
rect 55380 118880 55620 118900
rect 55880 118880 56120 118900
rect 56380 118880 56620 118900
rect 56880 118880 57120 118900
rect 57380 118880 57620 118900
rect 57880 118880 58000 118900
rect 14000 118620 14100 118880
rect 14400 118620 14600 118880
rect 14900 118620 15100 118880
rect 15400 118620 15600 118880
rect 15900 118620 16100 118880
rect 16400 118620 16600 118880
rect 16900 118620 17100 118880
rect 17400 118620 17600 118880
rect 17900 118620 18100 118880
rect 18400 118620 18600 118880
rect 18900 118620 19100 118880
rect 19400 118620 19600 118880
rect 19900 118620 20100 118880
rect 20400 118620 20600 118880
rect 20900 118620 21100 118880
rect 21400 118620 21600 118880
rect 21900 118620 22100 118880
rect 22400 118620 22600 118880
rect 22900 118620 23100 118880
rect 23400 118620 23600 118880
rect 23900 118620 24100 118880
rect 24400 118620 24600 118880
rect 24900 118620 25100 118880
rect 25400 118620 25600 118880
rect 25900 118620 26100 118880
rect 26400 118620 26600 118880
rect 26900 118620 27100 118880
rect 27400 118620 27600 118880
rect 27900 118620 28100 118880
rect 28400 118620 28600 118880
rect 28900 118620 29100 118880
rect 29400 118620 29600 118880
rect 29900 118620 30100 118880
rect 30400 118620 30600 118880
rect 30900 118620 31100 118880
rect 31400 118620 31600 118880
rect 31900 118620 32100 118880
rect 32400 118620 32600 118880
rect 32900 118620 33100 118880
rect 33400 118620 33600 118880
rect 33900 118620 34100 118880
rect 34400 118620 34600 118880
rect 34900 118620 35100 118880
rect 35400 118620 35600 118880
rect 35900 118620 36100 118880
rect 36400 118620 36600 118880
rect 36900 118620 37100 118880
rect 37400 118620 37600 118880
rect 37900 118620 38100 118880
rect 38400 118620 38600 118880
rect 38900 118620 39100 118880
rect 39400 118620 39600 118880
rect 39900 118620 40100 118880
rect 40400 118620 40600 118880
rect 40900 118620 41100 118880
rect 41400 118620 41600 118880
rect 41900 118620 42100 118880
rect 42400 118620 42600 118880
rect 42900 118620 43100 118880
rect 43400 118620 43600 118880
rect 43900 118620 44100 118880
rect 44400 118620 44600 118880
rect 44900 118620 45100 118880
rect 45400 118620 45600 118880
rect 45900 118620 46100 118880
rect 46400 118620 46600 118880
rect 46900 118620 47100 118880
rect 47400 118620 47600 118880
rect 47900 118620 48100 118880
rect 48400 118620 48600 118880
rect 48900 118620 49100 118880
rect 49400 118620 49600 118880
rect 49900 118620 50100 118880
rect 50400 118620 50600 118880
rect 50900 118620 51100 118880
rect 51400 118620 51600 118880
rect 51900 118620 52100 118880
rect 52400 118620 52600 118880
rect 52900 118620 53100 118880
rect 53400 118620 53600 118880
rect 53900 118620 54100 118880
rect 54400 118620 54600 118880
rect 54900 118620 55100 118880
rect 55400 118620 55600 118880
rect 55900 118620 56100 118880
rect 56400 118620 56600 118880
rect 56900 118620 57100 118880
rect 57400 118620 57600 118880
rect 57900 118620 58000 118880
rect 14000 118600 14120 118620
rect 14380 118600 14620 118620
rect 14880 118600 15120 118620
rect 15380 118600 15620 118620
rect 15880 118600 16120 118620
rect 16380 118600 16620 118620
rect 16880 118600 17120 118620
rect 17380 118600 17620 118620
rect 17880 118600 18120 118620
rect 18380 118600 18620 118620
rect 18880 118600 19120 118620
rect 19380 118600 19620 118620
rect 19880 118600 20120 118620
rect 20380 118600 20620 118620
rect 20880 118600 21120 118620
rect 21380 118600 21620 118620
rect 21880 118600 22120 118620
rect 22380 118600 22620 118620
rect 22880 118600 23120 118620
rect 23380 118600 23620 118620
rect 23880 118600 24120 118620
rect 24380 118600 24620 118620
rect 24880 118600 25120 118620
rect 25380 118600 25620 118620
rect 25880 118600 26120 118620
rect 26380 118600 26620 118620
rect 26880 118600 27120 118620
rect 27380 118600 27620 118620
rect 27880 118600 28120 118620
rect 28380 118600 28620 118620
rect 28880 118600 29120 118620
rect 29380 118600 29620 118620
rect 29880 118600 30120 118620
rect 30380 118600 30620 118620
rect 30880 118600 31120 118620
rect 31380 118600 31620 118620
rect 31880 118600 32120 118620
rect 32380 118600 32620 118620
rect 32880 118600 33120 118620
rect 33380 118600 33620 118620
rect 33880 118600 34120 118620
rect 34380 118600 34620 118620
rect 34880 118600 35120 118620
rect 35380 118600 35620 118620
rect 35880 118600 36120 118620
rect 36380 118600 36620 118620
rect 36880 118600 37120 118620
rect 37380 118600 37620 118620
rect 37880 118600 38120 118620
rect 38380 118600 38620 118620
rect 38880 118600 39120 118620
rect 39380 118600 39620 118620
rect 39880 118600 40120 118620
rect 40380 118600 40620 118620
rect 40880 118600 41120 118620
rect 41380 118600 41620 118620
rect 41880 118600 42120 118620
rect 42380 118600 42620 118620
rect 42880 118600 43120 118620
rect 43380 118600 43620 118620
rect 43880 118600 44120 118620
rect 44380 118600 44620 118620
rect 44880 118600 45120 118620
rect 45380 118600 45620 118620
rect 45880 118600 46120 118620
rect 46380 118600 46620 118620
rect 46880 118600 47120 118620
rect 47380 118600 47620 118620
rect 47880 118600 48120 118620
rect 48380 118600 48620 118620
rect 48880 118600 49120 118620
rect 49380 118600 49620 118620
rect 49880 118600 50120 118620
rect 50380 118600 50620 118620
rect 50880 118600 51120 118620
rect 51380 118600 51620 118620
rect 51880 118600 52120 118620
rect 52380 118600 52620 118620
rect 52880 118600 53120 118620
rect 53380 118600 53620 118620
rect 53880 118600 54120 118620
rect 54380 118600 54620 118620
rect 54880 118600 55120 118620
rect 55380 118600 55620 118620
rect 55880 118600 56120 118620
rect 56380 118600 56620 118620
rect 56880 118600 57120 118620
rect 57380 118600 57620 118620
rect 57880 118600 58000 118620
rect 14000 118400 58000 118600
rect 14000 118380 14120 118400
rect 14380 118380 14620 118400
rect 14880 118380 15120 118400
rect 15380 118380 15620 118400
rect 15880 118380 16120 118400
rect 16380 118380 16620 118400
rect 16880 118380 17120 118400
rect 17380 118380 17620 118400
rect 17880 118380 18120 118400
rect 18380 118380 18620 118400
rect 18880 118380 19120 118400
rect 19380 118380 19620 118400
rect 19880 118380 20120 118400
rect 20380 118380 20620 118400
rect 20880 118380 21120 118400
rect 21380 118380 21620 118400
rect 21880 118380 22120 118400
rect 22380 118380 22620 118400
rect 22880 118380 23120 118400
rect 23380 118380 23620 118400
rect 23880 118380 24120 118400
rect 24380 118380 24620 118400
rect 24880 118380 25120 118400
rect 25380 118380 25620 118400
rect 25880 118380 26120 118400
rect 26380 118380 26620 118400
rect 26880 118380 27120 118400
rect 27380 118380 27620 118400
rect 27880 118380 28120 118400
rect 28380 118380 28620 118400
rect 28880 118380 29120 118400
rect 29380 118380 29620 118400
rect 29880 118380 30120 118400
rect 30380 118380 30620 118400
rect 30880 118380 31120 118400
rect 31380 118380 31620 118400
rect 31880 118380 32120 118400
rect 32380 118380 32620 118400
rect 32880 118380 33120 118400
rect 33380 118380 33620 118400
rect 33880 118380 34120 118400
rect 34380 118380 34620 118400
rect 34880 118380 35120 118400
rect 35380 118380 35620 118400
rect 35880 118380 36120 118400
rect 36380 118380 36620 118400
rect 36880 118380 37120 118400
rect 37380 118380 37620 118400
rect 37880 118380 38120 118400
rect 38380 118380 38620 118400
rect 38880 118380 39120 118400
rect 39380 118380 39620 118400
rect 39880 118380 40120 118400
rect 40380 118380 40620 118400
rect 40880 118380 41120 118400
rect 41380 118380 41620 118400
rect 41880 118380 42120 118400
rect 42380 118380 42620 118400
rect 42880 118380 43120 118400
rect 43380 118380 43620 118400
rect 43880 118380 44120 118400
rect 44380 118380 44620 118400
rect 44880 118380 45120 118400
rect 45380 118380 45620 118400
rect 45880 118380 46120 118400
rect 46380 118380 46620 118400
rect 46880 118380 47120 118400
rect 47380 118380 47620 118400
rect 47880 118380 48120 118400
rect 48380 118380 48620 118400
rect 48880 118380 49120 118400
rect 49380 118380 49620 118400
rect 49880 118380 50120 118400
rect 50380 118380 50620 118400
rect 50880 118380 51120 118400
rect 51380 118380 51620 118400
rect 51880 118380 52120 118400
rect 52380 118380 52620 118400
rect 52880 118380 53120 118400
rect 53380 118380 53620 118400
rect 53880 118380 54120 118400
rect 54380 118380 54620 118400
rect 54880 118380 55120 118400
rect 55380 118380 55620 118400
rect 55880 118380 56120 118400
rect 56380 118380 56620 118400
rect 56880 118380 57120 118400
rect 57380 118380 57620 118400
rect 57880 118380 58000 118400
rect 14000 118120 14100 118380
rect 14400 118120 14600 118380
rect 14900 118120 15100 118380
rect 15400 118120 15600 118380
rect 15900 118120 16100 118380
rect 16400 118120 16600 118380
rect 16900 118120 17100 118380
rect 17400 118120 17600 118380
rect 17900 118120 18100 118380
rect 18400 118120 18600 118380
rect 18900 118120 19100 118380
rect 19400 118120 19600 118380
rect 19900 118120 20100 118380
rect 20400 118120 20600 118380
rect 20900 118120 21100 118380
rect 21400 118120 21600 118380
rect 21900 118120 22100 118380
rect 22400 118120 22600 118380
rect 22900 118120 23100 118380
rect 23400 118120 23600 118380
rect 23900 118120 24100 118380
rect 24400 118120 24600 118380
rect 24900 118120 25100 118380
rect 25400 118120 25600 118380
rect 25900 118120 26100 118380
rect 26400 118120 26600 118380
rect 26900 118120 27100 118380
rect 27400 118120 27600 118380
rect 27900 118120 28100 118380
rect 28400 118120 28600 118380
rect 28900 118120 29100 118380
rect 29400 118120 29600 118380
rect 29900 118120 30100 118380
rect 30400 118120 30600 118380
rect 30900 118120 31100 118380
rect 31400 118120 31600 118380
rect 31900 118120 32100 118380
rect 32400 118120 32600 118380
rect 32900 118120 33100 118380
rect 33400 118120 33600 118380
rect 33900 118120 34100 118380
rect 34400 118120 34600 118380
rect 34900 118120 35100 118380
rect 35400 118120 35600 118380
rect 35900 118120 36100 118380
rect 36400 118120 36600 118380
rect 36900 118120 37100 118380
rect 37400 118120 37600 118380
rect 37900 118120 38100 118380
rect 38400 118120 38600 118380
rect 38900 118120 39100 118380
rect 39400 118120 39600 118380
rect 39900 118120 40100 118380
rect 40400 118120 40600 118380
rect 40900 118120 41100 118380
rect 41400 118120 41600 118380
rect 41900 118120 42100 118380
rect 42400 118120 42600 118380
rect 42900 118120 43100 118380
rect 43400 118120 43600 118380
rect 43900 118120 44100 118380
rect 44400 118120 44600 118380
rect 44900 118120 45100 118380
rect 45400 118120 45600 118380
rect 45900 118120 46100 118380
rect 46400 118120 46600 118380
rect 46900 118120 47100 118380
rect 47400 118120 47600 118380
rect 47900 118120 48100 118380
rect 48400 118120 48600 118380
rect 48900 118120 49100 118380
rect 49400 118120 49600 118380
rect 49900 118120 50100 118380
rect 50400 118120 50600 118380
rect 50900 118120 51100 118380
rect 51400 118120 51600 118380
rect 51900 118120 52100 118380
rect 52400 118120 52600 118380
rect 52900 118120 53100 118380
rect 53400 118120 53600 118380
rect 53900 118120 54100 118380
rect 54400 118120 54600 118380
rect 54900 118120 55100 118380
rect 55400 118120 55600 118380
rect 55900 118120 56100 118380
rect 56400 118120 56600 118380
rect 56900 118120 57100 118380
rect 57400 118120 57600 118380
rect 57900 118120 58000 118380
rect 14000 118100 14120 118120
rect 14380 118100 14620 118120
rect 14880 118100 15120 118120
rect 15380 118100 15620 118120
rect 15880 118100 16120 118120
rect 16380 118100 16620 118120
rect 16880 118100 17120 118120
rect 17380 118100 17620 118120
rect 17880 118100 18120 118120
rect 18380 118100 18620 118120
rect 18880 118100 19120 118120
rect 19380 118100 19620 118120
rect 19880 118100 20120 118120
rect 20380 118100 20620 118120
rect 20880 118100 21120 118120
rect 21380 118100 21620 118120
rect 21880 118100 22120 118120
rect 22380 118100 22620 118120
rect 22880 118100 23120 118120
rect 23380 118100 23620 118120
rect 23880 118100 24120 118120
rect 24380 118100 24620 118120
rect 24880 118100 25120 118120
rect 25380 118100 25620 118120
rect 25880 118100 26120 118120
rect 26380 118100 26620 118120
rect 26880 118100 27120 118120
rect 27380 118100 27620 118120
rect 27880 118100 28120 118120
rect 28380 118100 28620 118120
rect 28880 118100 29120 118120
rect 29380 118100 29620 118120
rect 29880 118100 30120 118120
rect 30380 118100 30620 118120
rect 30880 118100 31120 118120
rect 31380 118100 31620 118120
rect 31880 118100 32120 118120
rect 32380 118100 32620 118120
rect 32880 118100 33120 118120
rect 33380 118100 33620 118120
rect 33880 118100 34120 118120
rect 34380 118100 34620 118120
rect 34880 118100 35120 118120
rect 35380 118100 35620 118120
rect 35880 118100 36120 118120
rect 36380 118100 36620 118120
rect 36880 118100 37120 118120
rect 37380 118100 37620 118120
rect 37880 118100 38120 118120
rect 38380 118100 38620 118120
rect 38880 118100 39120 118120
rect 39380 118100 39620 118120
rect 39880 118100 40120 118120
rect 40380 118100 40620 118120
rect 40880 118100 41120 118120
rect 41380 118100 41620 118120
rect 41880 118100 42120 118120
rect 42380 118100 42620 118120
rect 42880 118100 43120 118120
rect 43380 118100 43620 118120
rect 43880 118100 44120 118120
rect 44380 118100 44620 118120
rect 44880 118100 45120 118120
rect 45380 118100 45620 118120
rect 45880 118100 46120 118120
rect 46380 118100 46620 118120
rect 46880 118100 47120 118120
rect 47380 118100 47620 118120
rect 47880 118100 48120 118120
rect 48380 118100 48620 118120
rect 48880 118100 49120 118120
rect 49380 118100 49620 118120
rect 49880 118100 50120 118120
rect 50380 118100 50620 118120
rect 50880 118100 51120 118120
rect 51380 118100 51620 118120
rect 51880 118100 52120 118120
rect 52380 118100 52620 118120
rect 52880 118100 53120 118120
rect 53380 118100 53620 118120
rect 53880 118100 54120 118120
rect 54380 118100 54620 118120
rect 54880 118100 55120 118120
rect 55380 118100 55620 118120
rect 55880 118100 56120 118120
rect 56380 118100 56620 118120
rect 56880 118100 57120 118120
rect 57380 118100 57620 118120
rect 57880 118100 58000 118120
rect 14000 117900 58000 118100
rect 14000 117880 14120 117900
rect 14380 117880 14620 117900
rect 14880 117880 15120 117900
rect 15380 117880 15620 117900
rect 15880 117880 16120 117900
rect 16380 117880 16620 117900
rect 16880 117880 17120 117900
rect 17380 117880 17620 117900
rect 17880 117880 18120 117900
rect 18380 117880 18620 117900
rect 18880 117880 19120 117900
rect 19380 117880 19620 117900
rect 19880 117880 20120 117900
rect 20380 117880 20620 117900
rect 20880 117880 21120 117900
rect 21380 117880 21620 117900
rect 21880 117880 22120 117900
rect 22380 117880 22620 117900
rect 22880 117880 23120 117900
rect 23380 117880 23620 117900
rect 23880 117880 24120 117900
rect 24380 117880 24620 117900
rect 24880 117880 25120 117900
rect 25380 117880 25620 117900
rect 25880 117880 26120 117900
rect 26380 117880 26620 117900
rect 26880 117880 27120 117900
rect 27380 117880 27620 117900
rect 27880 117880 28120 117900
rect 28380 117880 28620 117900
rect 28880 117880 29120 117900
rect 29380 117880 29620 117900
rect 29880 117880 30120 117900
rect 30380 117880 30620 117900
rect 30880 117880 31120 117900
rect 31380 117880 31620 117900
rect 31880 117880 32120 117900
rect 32380 117880 32620 117900
rect 32880 117880 33120 117900
rect 33380 117880 33620 117900
rect 33880 117880 34120 117900
rect 34380 117880 34620 117900
rect 34880 117880 35120 117900
rect 35380 117880 35620 117900
rect 35880 117880 36120 117900
rect 36380 117880 36620 117900
rect 36880 117880 37120 117900
rect 37380 117880 37620 117900
rect 37880 117880 38120 117900
rect 38380 117880 38620 117900
rect 38880 117880 39120 117900
rect 39380 117880 39620 117900
rect 39880 117880 40120 117900
rect 40380 117880 40620 117900
rect 40880 117880 41120 117900
rect 41380 117880 41620 117900
rect 41880 117880 42120 117900
rect 42380 117880 42620 117900
rect 42880 117880 43120 117900
rect 43380 117880 43620 117900
rect 43880 117880 44120 117900
rect 44380 117880 44620 117900
rect 44880 117880 45120 117900
rect 45380 117880 45620 117900
rect 45880 117880 46120 117900
rect 46380 117880 46620 117900
rect 46880 117880 47120 117900
rect 47380 117880 47620 117900
rect 47880 117880 48120 117900
rect 48380 117880 48620 117900
rect 48880 117880 49120 117900
rect 49380 117880 49620 117900
rect 49880 117880 50120 117900
rect 50380 117880 50620 117900
rect 50880 117880 51120 117900
rect 51380 117880 51620 117900
rect 51880 117880 52120 117900
rect 52380 117880 52620 117900
rect 52880 117880 53120 117900
rect 53380 117880 53620 117900
rect 53880 117880 54120 117900
rect 54380 117880 54620 117900
rect 54880 117880 55120 117900
rect 55380 117880 55620 117900
rect 55880 117880 56120 117900
rect 56380 117880 56620 117900
rect 56880 117880 57120 117900
rect 57380 117880 57620 117900
rect 57880 117880 58000 117900
rect 14000 117620 14100 117880
rect 14400 117620 14600 117880
rect 14900 117620 15100 117880
rect 15400 117620 15600 117880
rect 15900 117620 16100 117880
rect 16400 117620 16600 117880
rect 16900 117620 17100 117880
rect 17400 117620 17600 117880
rect 17900 117620 18100 117880
rect 18400 117620 18600 117880
rect 18900 117620 19100 117880
rect 19400 117620 19600 117880
rect 19900 117620 20100 117880
rect 20400 117620 20600 117880
rect 20900 117620 21100 117880
rect 21400 117620 21600 117880
rect 21900 117620 22100 117880
rect 22400 117620 22600 117880
rect 22900 117620 23100 117880
rect 23400 117620 23600 117880
rect 23900 117620 24100 117880
rect 24400 117620 24600 117880
rect 24900 117620 25100 117880
rect 25400 117620 25600 117880
rect 25900 117620 26100 117880
rect 26400 117620 26600 117880
rect 26900 117620 27100 117880
rect 27400 117620 27600 117880
rect 27900 117620 28100 117880
rect 28400 117620 28600 117880
rect 28900 117620 29100 117880
rect 29400 117620 29600 117880
rect 29900 117620 30100 117880
rect 30400 117620 30600 117880
rect 30900 117620 31100 117880
rect 31400 117620 31600 117880
rect 31900 117620 32100 117880
rect 32400 117620 32600 117880
rect 32900 117620 33100 117880
rect 33400 117620 33600 117880
rect 33900 117620 34100 117880
rect 34400 117620 34600 117880
rect 34900 117620 35100 117880
rect 35400 117620 35600 117880
rect 35900 117620 36100 117880
rect 36400 117620 36600 117880
rect 36900 117620 37100 117880
rect 37400 117620 37600 117880
rect 37900 117620 38100 117880
rect 38400 117620 38600 117880
rect 38900 117620 39100 117880
rect 39400 117620 39600 117880
rect 39900 117620 40100 117880
rect 40400 117620 40600 117880
rect 40900 117620 41100 117880
rect 41400 117620 41600 117880
rect 41900 117620 42100 117880
rect 42400 117620 42600 117880
rect 42900 117620 43100 117880
rect 43400 117620 43600 117880
rect 43900 117620 44100 117880
rect 44400 117620 44600 117880
rect 44900 117620 45100 117880
rect 45400 117620 45600 117880
rect 45900 117620 46100 117880
rect 46400 117620 46600 117880
rect 46900 117620 47100 117880
rect 47400 117620 47600 117880
rect 47900 117620 48100 117880
rect 48400 117620 48600 117880
rect 48900 117620 49100 117880
rect 49400 117620 49600 117880
rect 49900 117620 50100 117880
rect 50400 117620 50600 117880
rect 50900 117620 51100 117880
rect 51400 117620 51600 117880
rect 51900 117620 52100 117880
rect 52400 117620 52600 117880
rect 52900 117620 53100 117880
rect 53400 117620 53600 117880
rect 53900 117620 54100 117880
rect 54400 117620 54600 117880
rect 54900 117620 55100 117880
rect 55400 117620 55600 117880
rect 55900 117620 56100 117880
rect 56400 117620 56600 117880
rect 56900 117620 57100 117880
rect 57400 117620 57600 117880
rect 57900 117620 58000 117880
rect 14000 117600 14120 117620
rect 14380 117600 14620 117620
rect 14880 117600 15120 117620
rect 15380 117600 15620 117620
rect 15880 117600 16120 117620
rect 16380 117600 16620 117620
rect 16880 117600 17120 117620
rect 17380 117600 17620 117620
rect 17880 117600 18120 117620
rect 18380 117600 18620 117620
rect 18880 117600 19120 117620
rect 19380 117600 19620 117620
rect 19880 117600 20120 117620
rect 20380 117600 20620 117620
rect 20880 117600 21120 117620
rect 21380 117600 21620 117620
rect 21880 117600 22120 117620
rect 22380 117600 22620 117620
rect 22880 117600 23120 117620
rect 23380 117600 23620 117620
rect 23880 117600 24120 117620
rect 24380 117600 24620 117620
rect 24880 117600 25120 117620
rect 25380 117600 25620 117620
rect 25880 117600 26120 117620
rect 26380 117600 26620 117620
rect 26880 117600 27120 117620
rect 27380 117600 27620 117620
rect 27880 117600 28120 117620
rect 28380 117600 28620 117620
rect 28880 117600 29120 117620
rect 29380 117600 29620 117620
rect 29880 117600 30120 117620
rect 30380 117600 30620 117620
rect 30880 117600 31120 117620
rect 31380 117600 31620 117620
rect 31880 117600 32120 117620
rect 32380 117600 32620 117620
rect 32880 117600 33120 117620
rect 33380 117600 33620 117620
rect 33880 117600 34120 117620
rect 34380 117600 34620 117620
rect 34880 117600 35120 117620
rect 35380 117600 35620 117620
rect 35880 117600 36120 117620
rect 36380 117600 36620 117620
rect 36880 117600 37120 117620
rect 37380 117600 37620 117620
rect 37880 117600 38120 117620
rect 38380 117600 38620 117620
rect 38880 117600 39120 117620
rect 39380 117600 39620 117620
rect 39880 117600 40120 117620
rect 40380 117600 40620 117620
rect 40880 117600 41120 117620
rect 41380 117600 41620 117620
rect 41880 117600 42120 117620
rect 42380 117600 42620 117620
rect 42880 117600 43120 117620
rect 43380 117600 43620 117620
rect 43880 117600 44120 117620
rect 44380 117600 44620 117620
rect 44880 117600 45120 117620
rect 45380 117600 45620 117620
rect 45880 117600 46120 117620
rect 46380 117600 46620 117620
rect 46880 117600 47120 117620
rect 47380 117600 47620 117620
rect 47880 117600 48120 117620
rect 48380 117600 48620 117620
rect 48880 117600 49120 117620
rect 49380 117600 49620 117620
rect 49880 117600 50120 117620
rect 50380 117600 50620 117620
rect 50880 117600 51120 117620
rect 51380 117600 51620 117620
rect 51880 117600 52120 117620
rect 52380 117600 52620 117620
rect 52880 117600 53120 117620
rect 53380 117600 53620 117620
rect 53880 117600 54120 117620
rect 54380 117600 54620 117620
rect 54880 117600 55120 117620
rect 55380 117600 55620 117620
rect 55880 117600 56120 117620
rect 56380 117600 56620 117620
rect 56880 117600 57120 117620
rect 57380 117600 57620 117620
rect 57880 117600 58000 117620
rect 14000 117400 58000 117600
rect 14000 117380 14120 117400
rect 14380 117380 14620 117400
rect 14880 117380 15120 117400
rect 15380 117380 15620 117400
rect 15880 117380 16120 117400
rect 16380 117380 16620 117400
rect 16880 117380 17120 117400
rect 17380 117380 17620 117400
rect 17880 117380 18120 117400
rect 18380 117380 18620 117400
rect 18880 117380 19120 117400
rect 19380 117380 19620 117400
rect 19880 117380 20120 117400
rect 20380 117380 20620 117400
rect 20880 117380 21120 117400
rect 21380 117380 21620 117400
rect 21880 117380 22120 117400
rect 22380 117380 22620 117400
rect 22880 117380 23120 117400
rect 23380 117380 23620 117400
rect 23880 117380 24120 117400
rect 24380 117380 24620 117400
rect 24880 117380 25120 117400
rect 25380 117380 25620 117400
rect 25880 117380 26120 117400
rect 26380 117380 26620 117400
rect 26880 117380 27120 117400
rect 27380 117380 27620 117400
rect 27880 117380 28120 117400
rect 28380 117380 28620 117400
rect 28880 117380 29120 117400
rect 29380 117380 29620 117400
rect 29880 117380 30120 117400
rect 30380 117380 30620 117400
rect 30880 117380 31120 117400
rect 31380 117380 31620 117400
rect 31880 117380 32120 117400
rect 32380 117380 32620 117400
rect 32880 117380 33120 117400
rect 33380 117380 33620 117400
rect 33880 117380 34120 117400
rect 34380 117380 34620 117400
rect 34880 117380 35120 117400
rect 35380 117380 35620 117400
rect 35880 117380 36120 117400
rect 36380 117380 36620 117400
rect 36880 117380 37120 117400
rect 37380 117380 37620 117400
rect 37880 117380 38120 117400
rect 38380 117380 38620 117400
rect 38880 117380 39120 117400
rect 39380 117380 39620 117400
rect 39880 117380 40120 117400
rect 40380 117380 40620 117400
rect 40880 117380 41120 117400
rect 41380 117380 41620 117400
rect 41880 117380 42120 117400
rect 42380 117380 42620 117400
rect 42880 117380 43120 117400
rect 43380 117380 43620 117400
rect 43880 117380 44120 117400
rect 44380 117380 44620 117400
rect 44880 117380 45120 117400
rect 45380 117380 45620 117400
rect 45880 117380 46120 117400
rect 46380 117380 46620 117400
rect 46880 117380 47120 117400
rect 47380 117380 47620 117400
rect 47880 117380 48120 117400
rect 48380 117380 48620 117400
rect 48880 117380 49120 117400
rect 49380 117380 49620 117400
rect 49880 117380 50120 117400
rect 50380 117380 50620 117400
rect 50880 117380 51120 117400
rect 51380 117380 51620 117400
rect 51880 117380 52120 117400
rect 52380 117380 52620 117400
rect 52880 117380 53120 117400
rect 53380 117380 53620 117400
rect 53880 117380 54120 117400
rect 54380 117380 54620 117400
rect 54880 117380 55120 117400
rect 55380 117380 55620 117400
rect 55880 117380 56120 117400
rect 56380 117380 56620 117400
rect 56880 117380 57120 117400
rect 57380 117380 57620 117400
rect 57880 117380 58000 117400
rect 14000 117120 14100 117380
rect 14400 117120 14600 117380
rect 14900 117120 15100 117380
rect 15400 117120 15600 117380
rect 15900 117120 16100 117380
rect 16400 117120 16600 117380
rect 16900 117120 17100 117380
rect 17400 117120 17600 117380
rect 17900 117120 18100 117380
rect 18400 117120 18600 117380
rect 18900 117120 19100 117380
rect 19400 117120 19600 117380
rect 19900 117120 20100 117380
rect 20400 117120 20600 117380
rect 20900 117120 21100 117380
rect 21400 117120 21600 117380
rect 21900 117120 22100 117380
rect 22400 117120 22600 117380
rect 22900 117120 23100 117380
rect 23400 117120 23600 117380
rect 23900 117120 24100 117380
rect 24400 117120 24600 117380
rect 24900 117120 25100 117380
rect 25400 117120 25600 117380
rect 25900 117120 26100 117380
rect 26400 117120 26600 117380
rect 26900 117120 27100 117380
rect 27400 117120 27600 117380
rect 27900 117120 28100 117380
rect 28400 117120 28600 117380
rect 28900 117120 29100 117380
rect 29400 117120 29600 117380
rect 29900 117120 30100 117380
rect 30400 117120 30600 117380
rect 30900 117120 31100 117380
rect 31400 117120 31600 117380
rect 31900 117120 32100 117380
rect 32400 117120 32600 117380
rect 32900 117120 33100 117380
rect 33400 117120 33600 117380
rect 33900 117120 34100 117380
rect 34400 117120 34600 117380
rect 34900 117120 35100 117380
rect 35400 117120 35600 117380
rect 35900 117120 36100 117380
rect 36400 117120 36600 117380
rect 36900 117120 37100 117380
rect 37400 117120 37600 117380
rect 37900 117120 38100 117380
rect 38400 117120 38600 117380
rect 38900 117120 39100 117380
rect 39400 117120 39600 117380
rect 39900 117120 40100 117380
rect 40400 117120 40600 117380
rect 40900 117120 41100 117380
rect 41400 117120 41600 117380
rect 41900 117120 42100 117380
rect 42400 117120 42600 117380
rect 42900 117120 43100 117380
rect 43400 117120 43600 117380
rect 43900 117120 44100 117380
rect 44400 117120 44600 117380
rect 44900 117120 45100 117380
rect 45400 117120 45600 117380
rect 45900 117120 46100 117380
rect 46400 117120 46600 117380
rect 46900 117120 47100 117380
rect 47400 117120 47600 117380
rect 47900 117120 48100 117380
rect 48400 117120 48600 117380
rect 48900 117120 49100 117380
rect 49400 117120 49600 117380
rect 49900 117120 50100 117380
rect 50400 117120 50600 117380
rect 50900 117120 51100 117380
rect 51400 117120 51600 117380
rect 51900 117120 52100 117380
rect 52400 117120 52600 117380
rect 52900 117120 53100 117380
rect 53400 117120 53600 117380
rect 53900 117120 54100 117380
rect 54400 117120 54600 117380
rect 54900 117120 55100 117380
rect 55400 117120 55600 117380
rect 55900 117120 56100 117380
rect 56400 117120 56600 117380
rect 56900 117120 57100 117380
rect 57400 117120 57600 117380
rect 57900 117120 58000 117380
rect 14000 117100 14120 117120
rect 14380 117100 14620 117120
rect 14880 117100 15120 117120
rect 15380 117100 15620 117120
rect 15880 117100 16120 117120
rect 16380 117100 16620 117120
rect 16880 117100 17120 117120
rect 17380 117100 17620 117120
rect 17880 117100 18120 117120
rect 18380 117100 18620 117120
rect 18880 117100 19120 117120
rect 19380 117100 19620 117120
rect 19880 117100 20120 117120
rect 20380 117100 20620 117120
rect 20880 117100 21120 117120
rect 21380 117100 21620 117120
rect 21880 117100 22120 117120
rect 22380 117100 22620 117120
rect 22880 117100 23120 117120
rect 23380 117100 23620 117120
rect 23880 117100 24120 117120
rect 24380 117100 24620 117120
rect 24880 117100 25120 117120
rect 25380 117100 25620 117120
rect 25880 117100 26120 117120
rect 26380 117100 26620 117120
rect 26880 117100 27120 117120
rect 27380 117100 27620 117120
rect 27880 117100 28120 117120
rect 28380 117100 28620 117120
rect 28880 117100 29120 117120
rect 29380 117100 29620 117120
rect 29880 117100 30120 117120
rect 30380 117100 30620 117120
rect 30880 117100 31120 117120
rect 31380 117100 31620 117120
rect 31880 117100 32120 117120
rect 32380 117100 32620 117120
rect 32880 117100 33120 117120
rect 33380 117100 33620 117120
rect 33880 117100 34120 117120
rect 34380 117100 34620 117120
rect 34880 117100 35120 117120
rect 35380 117100 35620 117120
rect 35880 117100 36120 117120
rect 36380 117100 36620 117120
rect 36880 117100 37120 117120
rect 37380 117100 37620 117120
rect 37880 117100 38120 117120
rect 38380 117100 38620 117120
rect 38880 117100 39120 117120
rect 39380 117100 39620 117120
rect 39880 117100 40120 117120
rect 40380 117100 40620 117120
rect 40880 117100 41120 117120
rect 41380 117100 41620 117120
rect 41880 117100 42120 117120
rect 42380 117100 42620 117120
rect 42880 117100 43120 117120
rect 43380 117100 43620 117120
rect 43880 117100 44120 117120
rect 44380 117100 44620 117120
rect 44880 117100 45120 117120
rect 45380 117100 45620 117120
rect 45880 117100 46120 117120
rect 46380 117100 46620 117120
rect 46880 117100 47120 117120
rect 47380 117100 47620 117120
rect 47880 117100 48120 117120
rect 48380 117100 48620 117120
rect 48880 117100 49120 117120
rect 49380 117100 49620 117120
rect 49880 117100 50120 117120
rect 50380 117100 50620 117120
rect 50880 117100 51120 117120
rect 51380 117100 51620 117120
rect 51880 117100 52120 117120
rect 52380 117100 52620 117120
rect 52880 117100 53120 117120
rect 53380 117100 53620 117120
rect 53880 117100 54120 117120
rect 54380 117100 54620 117120
rect 54880 117100 55120 117120
rect 55380 117100 55620 117120
rect 55880 117100 56120 117120
rect 56380 117100 56620 117120
rect 56880 117100 57120 117120
rect 57380 117100 57620 117120
rect 57880 117100 58000 117120
rect 14000 116900 58000 117100
rect 14000 116880 14120 116900
rect 14380 116880 14620 116900
rect 14880 116880 15120 116900
rect 15380 116880 15620 116900
rect 15880 116880 16120 116900
rect 16380 116880 16620 116900
rect 16880 116880 17120 116900
rect 17380 116880 17620 116900
rect 17880 116880 18120 116900
rect 18380 116880 18620 116900
rect 18880 116880 19120 116900
rect 19380 116880 19620 116900
rect 19880 116880 20120 116900
rect 20380 116880 20620 116900
rect 20880 116880 21120 116900
rect 21380 116880 21620 116900
rect 21880 116880 22120 116900
rect 22380 116880 22620 116900
rect 22880 116880 23120 116900
rect 23380 116880 23620 116900
rect 23880 116880 24120 116900
rect 24380 116880 24620 116900
rect 24880 116880 25120 116900
rect 25380 116880 25620 116900
rect 25880 116880 26120 116900
rect 26380 116880 26620 116900
rect 26880 116880 27120 116900
rect 27380 116880 27620 116900
rect 27880 116880 28120 116900
rect 28380 116880 28620 116900
rect 28880 116880 29120 116900
rect 29380 116880 29620 116900
rect 29880 116880 30120 116900
rect 30380 116880 30620 116900
rect 30880 116880 31120 116900
rect 31380 116880 31620 116900
rect 31880 116880 32120 116900
rect 32380 116880 32620 116900
rect 32880 116880 33120 116900
rect 33380 116880 33620 116900
rect 33880 116880 34120 116900
rect 34380 116880 34620 116900
rect 34880 116880 35120 116900
rect 35380 116880 35620 116900
rect 35880 116880 36120 116900
rect 36380 116880 36620 116900
rect 36880 116880 37120 116900
rect 37380 116880 37620 116900
rect 37880 116880 38120 116900
rect 38380 116880 38620 116900
rect 38880 116880 39120 116900
rect 39380 116880 39620 116900
rect 39880 116880 40120 116900
rect 40380 116880 40620 116900
rect 40880 116880 41120 116900
rect 41380 116880 41620 116900
rect 41880 116880 42120 116900
rect 42380 116880 42620 116900
rect 42880 116880 43120 116900
rect 43380 116880 43620 116900
rect 43880 116880 44120 116900
rect 44380 116880 44620 116900
rect 44880 116880 45120 116900
rect 45380 116880 45620 116900
rect 45880 116880 46120 116900
rect 46380 116880 46620 116900
rect 46880 116880 47120 116900
rect 47380 116880 47620 116900
rect 47880 116880 48120 116900
rect 48380 116880 48620 116900
rect 48880 116880 49120 116900
rect 49380 116880 49620 116900
rect 49880 116880 50120 116900
rect 50380 116880 50620 116900
rect 50880 116880 51120 116900
rect 51380 116880 51620 116900
rect 51880 116880 52120 116900
rect 52380 116880 52620 116900
rect 52880 116880 53120 116900
rect 53380 116880 53620 116900
rect 53880 116880 54120 116900
rect 54380 116880 54620 116900
rect 54880 116880 55120 116900
rect 55380 116880 55620 116900
rect 55880 116880 56120 116900
rect 56380 116880 56620 116900
rect 56880 116880 57120 116900
rect 57380 116880 57620 116900
rect 57880 116880 58000 116900
rect 14000 116620 14100 116880
rect 14400 116620 14600 116880
rect 14900 116620 15100 116880
rect 15400 116620 15600 116880
rect 15900 116620 16100 116880
rect 16400 116620 16600 116880
rect 16900 116620 17100 116880
rect 17400 116620 17600 116880
rect 17900 116620 18100 116880
rect 18400 116620 18600 116880
rect 18900 116620 19100 116880
rect 19400 116620 19600 116880
rect 19900 116620 20100 116880
rect 20400 116620 20600 116880
rect 20900 116620 21100 116880
rect 21400 116620 21600 116880
rect 21900 116620 22100 116880
rect 22400 116620 22600 116880
rect 22900 116620 23100 116880
rect 23400 116620 23600 116880
rect 23900 116620 24100 116880
rect 24400 116620 24600 116880
rect 24900 116620 25100 116880
rect 25400 116620 25600 116880
rect 25900 116620 26100 116880
rect 26400 116620 26600 116880
rect 26900 116620 27100 116880
rect 27400 116620 27600 116880
rect 27900 116620 28100 116880
rect 28400 116620 28600 116880
rect 28900 116620 29100 116880
rect 29400 116620 29600 116880
rect 29900 116620 30100 116880
rect 30400 116620 30600 116880
rect 30900 116620 31100 116880
rect 31400 116620 31600 116880
rect 31900 116620 32100 116880
rect 32400 116620 32600 116880
rect 32900 116620 33100 116880
rect 33400 116620 33600 116880
rect 33900 116620 34100 116880
rect 34400 116620 34600 116880
rect 34900 116620 35100 116880
rect 35400 116620 35600 116880
rect 35900 116620 36100 116880
rect 36400 116620 36600 116880
rect 36900 116620 37100 116880
rect 37400 116620 37600 116880
rect 37900 116620 38100 116880
rect 38400 116620 38600 116880
rect 38900 116620 39100 116880
rect 39400 116620 39600 116880
rect 39900 116620 40100 116880
rect 40400 116620 40600 116880
rect 40900 116620 41100 116880
rect 41400 116620 41600 116880
rect 41900 116620 42100 116880
rect 42400 116620 42600 116880
rect 42900 116620 43100 116880
rect 43400 116620 43600 116880
rect 43900 116620 44100 116880
rect 44400 116620 44600 116880
rect 44900 116620 45100 116880
rect 45400 116620 45600 116880
rect 45900 116620 46100 116880
rect 46400 116620 46600 116880
rect 46900 116620 47100 116880
rect 47400 116620 47600 116880
rect 47900 116620 48100 116880
rect 48400 116620 48600 116880
rect 48900 116620 49100 116880
rect 49400 116620 49600 116880
rect 49900 116620 50100 116880
rect 50400 116620 50600 116880
rect 50900 116620 51100 116880
rect 51400 116620 51600 116880
rect 51900 116620 52100 116880
rect 52400 116620 52600 116880
rect 52900 116620 53100 116880
rect 53400 116620 53600 116880
rect 53900 116620 54100 116880
rect 54400 116620 54600 116880
rect 54900 116620 55100 116880
rect 55400 116620 55600 116880
rect 55900 116620 56100 116880
rect 56400 116620 56600 116880
rect 56900 116620 57100 116880
rect 57400 116620 57600 116880
rect 57900 116620 58000 116880
rect 14000 116600 14120 116620
rect 14380 116600 14620 116620
rect 14880 116600 15120 116620
rect 15380 116600 15620 116620
rect 15880 116600 16120 116620
rect 16380 116600 16620 116620
rect 16880 116600 17120 116620
rect 17380 116600 17620 116620
rect 17880 116600 18120 116620
rect 18380 116600 18620 116620
rect 18880 116600 19120 116620
rect 19380 116600 19620 116620
rect 19880 116600 20120 116620
rect 20380 116600 20620 116620
rect 20880 116600 21120 116620
rect 21380 116600 21620 116620
rect 21880 116600 22120 116620
rect 22380 116600 22620 116620
rect 22880 116600 23120 116620
rect 23380 116600 23620 116620
rect 23880 116600 24120 116620
rect 24380 116600 24620 116620
rect 24880 116600 25120 116620
rect 25380 116600 25620 116620
rect 25880 116600 26120 116620
rect 26380 116600 26620 116620
rect 26880 116600 27120 116620
rect 27380 116600 27620 116620
rect 27880 116600 28120 116620
rect 28380 116600 28620 116620
rect 28880 116600 29120 116620
rect 29380 116600 29620 116620
rect 29880 116600 30120 116620
rect 30380 116600 30620 116620
rect 30880 116600 31120 116620
rect 31380 116600 31620 116620
rect 31880 116600 32120 116620
rect 32380 116600 32620 116620
rect 32880 116600 33120 116620
rect 33380 116600 33620 116620
rect 33880 116600 34120 116620
rect 34380 116600 34620 116620
rect 34880 116600 35120 116620
rect 35380 116600 35620 116620
rect 35880 116600 36120 116620
rect 36380 116600 36620 116620
rect 36880 116600 37120 116620
rect 37380 116600 37620 116620
rect 37880 116600 38120 116620
rect 38380 116600 38620 116620
rect 38880 116600 39120 116620
rect 39380 116600 39620 116620
rect 39880 116600 40120 116620
rect 40380 116600 40620 116620
rect 40880 116600 41120 116620
rect 41380 116600 41620 116620
rect 41880 116600 42120 116620
rect 42380 116600 42620 116620
rect 42880 116600 43120 116620
rect 43380 116600 43620 116620
rect 43880 116600 44120 116620
rect 44380 116600 44620 116620
rect 44880 116600 45120 116620
rect 45380 116600 45620 116620
rect 45880 116600 46120 116620
rect 46380 116600 46620 116620
rect 46880 116600 47120 116620
rect 47380 116600 47620 116620
rect 47880 116600 48120 116620
rect 48380 116600 48620 116620
rect 48880 116600 49120 116620
rect 49380 116600 49620 116620
rect 49880 116600 50120 116620
rect 50380 116600 50620 116620
rect 50880 116600 51120 116620
rect 51380 116600 51620 116620
rect 51880 116600 52120 116620
rect 52380 116600 52620 116620
rect 52880 116600 53120 116620
rect 53380 116600 53620 116620
rect 53880 116600 54120 116620
rect 54380 116600 54620 116620
rect 54880 116600 55120 116620
rect 55380 116600 55620 116620
rect 55880 116600 56120 116620
rect 56380 116600 56620 116620
rect 56880 116600 57120 116620
rect 57380 116600 57620 116620
rect 57880 116600 58000 116620
rect 14000 116400 58000 116600
rect 14000 116380 14120 116400
rect 14380 116380 14620 116400
rect 14880 116380 15120 116400
rect 15380 116380 15620 116400
rect 15880 116380 16120 116400
rect 16380 116380 16620 116400
rect 16880 116380 17120 116400
rect 17380 116380 17620 116400
rect 17880 116380 18120 116400
rect 18380 116380 18620 116400
rect 18880 116380 19120 116400
rect 19380 116380 19620 116400
rect 19880 116380 20120 116400
rect 20380 116380 20620 116400
rect 20880 116380 21120 116400
rect 21380 116380 21620 116400
rect 21880 116380 22120 116400
rect 22380 116380 22620 116400
rect 22880 116380 23120 116400
rect 23380 116380 23620 116400
rect 23880 116380 24120 116400
rect 24380 116380 24620 116400
rect 24880 116380 25120 116400
rect 25380 116380 25620 116400
rect 25880 116380 26120 116400
rect 26380 116380 26620 116400
rect 26880 116380 27120 116400
rect 27380 116380 27620 116400
rect 27880 116380 28120 116400
rect 28380 116380 28620 116400
rect 28880 116380 29120 116400
rect 29380 116380 29620 116400
rect 29880 116380 30120 116400
rect 30380 116380 30620 116400
rect 30880 116380 31120 116400
rect 31380 116380 31620 116400
rect 31880 116380 32120 116400
rect 32380 116380 32620 116400
rect 32880 116380 33120 116400
rect 33380 116380 33620 116400
rect 33880 116380 34120 116400
rect 34380 116380 34620 116400
rect 34880 116380 35120 116400
rect 35380 116380 35620 116400
rect 35880 116380 36120 116400
rect 36380 116380 36620 116400
rect 36880 116380 37120 116400
rect 37380 116380 37620 116400
rect 37880 116380 38120 116400
rect 38380 116380 38620 116400
rect 38880 116380 39120 116400
rect 39380 116380 39620 116400
rect 39880 116380 40120 116400
rect 40380 116380 40620 116400
rect 40880 116380 41120 116400
rect 41380 116380 41620 116400
rect 41880 116380 42120 116400
rect 42380 116380 42620 116400
rect 42880 116380 43120 116400
rect 43380 116380 43620 116400
rect 43880 116380 44120 116400
rect 44380 116380 44620 116400
rect 44880 116380 45120 116400
rect 45380 116380 45620 116400
rect 45880 116380 46120 116400
rect 46380 116380 46620 116400
rect 46880 116380 47120 116400
rect 47380 116380 47620 116400
rect 47880 116380 48120 116400
rect 48380 116380 48620 116400
rect 48880 116380 49120 116400
rect 49380 116380 49620 116400
rect 49880 116380 50120 116400
rect 50380 116380 50620 116400
rect 50880 116380 51120 116400
rect 51380 116380 51620 116400
rect 51880 116380 52120 116400
rect 52380 116380 52620 116400
rect 52880 116380 53120 116400
rect 53380 116380 53620 116400
rect 53880 116380 54120 116400
rect 54380 116380 54620 116400
rect 54880 116380 55120 116400
rect 55380 116380 55620 116400
rect 55880 116380 56120 116400
rect 56380 116380 56620 116400
rect 56880 116380 57120 116400
rect 57380 116380 57620 116400
rect 57880 116380 58000 116400
rect 14000 116120 14100 116380
rect 14400 116120 14600 116380
rect 14900 116120 15100 116380
rect 15400 116120 15600 116380
rect 15900 116120 16100 116380
rect 16400 116120 16600 116380
rect 16900 116120 17100 116380
rect 17400 116120 17600 116380
rect 17900 116120 18100 116380
rect 18400 116120 18600 116380
rect 18900 116120 19100 116380
rect 19400 116120 19600 116380
rect 19900 116120 20100 116380
rect 20400 116120 20600 116380
rect 20900 116120 21100 116380
rect 21400 116120 21600 116380
rect 21900 116120 22100 116380
rect 22400 116120 22600 116380
rect 22900 116120 23100 116380
rect 23400 116120 23600 116380
rect 23900 116120 24100 116380
rect 24400 116120 24600 116380
rect 24900 116120 25100 116380
rect 25400 116120 25600 116380
rect 25900 116120 26100 116380
rect 26400 116120 26600 116380
rect 26900 116120 27100 116380
rect 27400 116120 27600 116380
rect 27900 116120 28100 116380
rect 28400 116120 28600 116380
rect 28900 116120 29100 116380
rect 29400 116120 29600 116380
rect 29900 116120 30100 116380
rect 30400 116120 30600 116380
rect 30900 116120 31100 116380
rect 31400 116120 31600 116380
rect 31900 116120 32100 116380
rect 32400 116120 32600 116380
rect 32900 116120 33100 116380
rect 33400 116120 33600 116380
rect 33900 116120 34100 116380
rect 34400 116120 34600 116380
rect 34900 116120 35100 116380
rect 35400 116120 35600 116380
rect 35900 116120 36100 116380
rect 36400 116120 36600 116380
rect 36900 116120 37100 116380
rect 37400 116120 37600 116380
rect 37900 116120 38100 116380
rect 38400 116120 38600 116380
rect 38900 116120 39100 116380
rect 39400 116120 39600 116380
rect 39900 116120 40100 116380
rect 40400 116120 40600 116380
rect 40900 116120 41100 116380
rect 41400 116120 41600 116380
rect 41900 116120 42100 116380
rect 42400 116120 42600 116380
rect 42900 116120 43100 116380
rect 43400 116120 43600 116380
rect 43900 116120 44100 116380
rect 44400 116120 44600 116380
rect 44900 116120 45100 116380
rect 45400 116120 45600 116380
rect 45900 116120 46100 116380
rect 46400 116120 46600 116380
rect 46900 116120 47100 116380
rect 47400 116120 47600 116380
rect 47900 116120 48100 116380
rect 48400 116120 48600 116380
rect 48900 116120 49100 116380
rect 49400 116120 49600 116380
rect 49900 116120 50100 116380
rect 50400 116120 50600 116380
rect 50900 116120 51100 116380
rect 51400 116120 51600 116380
rect 51900 116120 52100 116380
rect 52400 116120 52600 116380
rect 52900 116120 53100 116380
rect 53400 116120 53600 116380
rect 53900 116120 54100 116380
rect 54400 116120 54600 116380
rect 54900 116120 55100 116380
rect 55400 116120 55600 116380
rect 55900 116120 56100 116380
rect 56400 116120 56600 116380
rect 56900 116120 57100 116380
rect 57400 116120 57600 116380
rect 57900 116120 58000 116380
rect 14000 116100 14120 116120
rect 14380 116100 14620 116120
rect 14880 116100 15120 116120
rect 15380 116100 15620 116120
rect 15880 116100 16120 116120
rect 16380 116100 16620 116120
rect 16880 116100 17120 116120
rect 17380 116100 17620 116120
rect 17880 116100 18120 116120
rect 18380 116100 18620 116120
rect 18880 116100 19120 116120
rect 19380 116100 19620 116120
rect 19880 116100 20120 116120
rect 20380 116100 20620 116120
rect 20880 116100 21120 116120
rect 21380 116100 21620 116120
rect 21880 116100 22120 116120
rect 22380 116100 22620 116120
rect 22880 116100 23120 116120
rect 23380 116100 23620 116120
rect 23880 116100 24120 116120
rect 24380 116100 24620 116120
rect 24880 116100 25120 116120
rect 25380 116100 25620 116120
rect 25880 116100 26120 116120
rect 26380 116100 26620 116120
rect 26880 116100 27120 116120
rect 27380 116100 27620 116120
rect 27880 116100 28120 116120
rect 28380 116100 28620 116120
rect 28880 116100 29120 116120
rect 29380 116100 29620 116120
rect 29880 116100 30120 116120
rect 30380 116100 30620 116120
rect 30880 116100 31120 116120
rect 31380 116100 31620 116120
rect 31880 116100 32120 116120
rect 32380 116100 32620 116120
rect 32880 116100 33120 116120
rect 33380 116100 33620 116120
rect 33880 116100 34120 116120
rect 34380 116100 34620 116120
rect 34880 116100 35120 116120
rect 35380 116100 35620 116120
rect 35880 116100 36120 116120
rect 36380 116100 36620 116120
rect 36880 116100 37120 116120
rect 37380 116100 37620 116120
rect 37880 116100 38120 116120
rect 38380 116100 38620 116120
rect 38880 116100 39120 116120
rect 39380 116100 39620 116120
rect 39880 116100 40120 116120
rect 40380 116100 40620 116120
rect 40880 116100 41120 116120
rect 41380 116100 41620 116120
rect 41880 116100 42120 116120
rect 42380 116100 42620 116120
rect 42880 116100 43120 116120
rect 43380 116100 43620 116120
rect 43880 116100 44120 116120
rect 44380 116100 44620 116120
rect 44880 116100 45120 116120
rect 45380 116100 45620 116120
rect 45880 116100 46120 116120
rect 46380 116100 46620 116120
rect 46880 116100 47120 116120
rect 47380 116100 47620 116120
rect 47880 116100 48120 116120
rect 48380 116100 48620 116120
rect 48880 116100 49120 116120
rect 49380 116100 49620 116120
rect 49880 116100 50120 116120
rect 50380 116100 50620 116120
rect 50880 116100 51120 116120
rect 51380 116100 51620 116120
rect 51880 116100 52120 116120
rect 52380 116100 52620 116120
rect 52880 116100 53120 116120
rect 53380 116100 53620 116120
rect 53880 116100 54120 116120
rect 54380 116100 54620 116120
rect 54880 116100 55120 116120
rect 55380 116100 55620 116120
rect 55880 116100 56120 116120
rect 56380 116100 56620 116120
rect 56880 116100 57120 116120
rect 57380 116100 57620 116120
rect 57880 116100 58000 116120
rect 14000 115900 58000 116100
rect 14000 115880 14120 115900
rect 14380 115880 14620 115900
rect 14880 115880 15120 115900
rect 15380 115880 15620 115900
rect 15880 115880 16120 115900
rect 16380 115880 16620 115900
rect 16880 115880 17120 115900
rect 17380 115880 17620 115900
rect 17880 115880 18120 115900
rect 18380 115880 18620 115900
rect 18880 115880 19120 115900
rect 19380 115880 19620 115900
rect 19880 115880 20120 115900
rect 20380 115880 20620 115900
rect 20880 115880 21120 115900
rect 21380 115880 21620 115900
rect 21880 115880 22120 115900
rect 22380 115880 22620 115900
rect 22880 115880 23120 115900
rect 23380 115880 23620 115900
rect 23880 115880 24120 115900
rect 24380 115880 24620 115900
rect 24880 115880 25120 115900
rect 25380 115880 25620 115900
rect 25880 115880 26120 115900
rect 26380 115880 26620 115900
rect 26880 115880 27120 115900
rect 27380 115880 27620 115900
rect 27880 115880 28120 115900
rect 28380 115880 28620 115900
rect 28880 115880 29120 115900
rect 29380 115880 29620 115900
rect 29880 115880 30120 115900
rect 30380 115880 30620 115900
rect 30880 115880 31120 115900
rect 31380 115880 31620 115900
rect 31880 115880 32120 115900
rect 32380 115880 32620 115900
rect 32880 115880 33120 115900
rect 33380 115880 33620 115900
rect 33880 115880 34120 115900
rect 34380 115880 34620 115900
rect 34880 115880 35120 115900
rect 35380 115880 35620 115900
rect 35880 115880 36120 115900
rect 36380 115880 36620 115900
rect 36880 115880 37120 115900
rect 37380 115880 37620 115900
rect 37880 115880 38120 115900
rect 38380 115880 38620 115900
rect 38880 115880 39120 115900
rect 39380 115880 39620 115900
rect 39880 115880 40120 115900
rect 40380 115880 40620 115900
rect 40880 115880 41120 115900
rect 41380 115880 41620 115900
rect 41880 115880 42120 115900
rect 42380 115880 42620 115900
rect 42880 115880 43120 115900
rect 43380 115880 43620 115900
rect 43880 115880 44120 115900
rect 44380 115880 44620 115900
rect 44880 115880 45120 115900
rect 45380 115880 45620 115900
rect 45880 115880 46120 115900
rect 46380 115880 46620 115900
rect 46880 115880 47120 115900
rect 47380 115880 47620 115900
rect 47880 115880 48120 115900
rect 48380 115880 48620 115900
rect 48880 115880 49120 115900
rect 49380 115880 49620 115900
rect 49880 115880 50120 115900
rect 50380 115880 50620 115900
rect 50880 115880 51120 115900
rect 51380 115880 51620 115900
rect 51880 115880 52120 115900
rect 52380 115880 52620 115900
rect 52880 115880 53120 115900
rect 53380 115880 53620 115900
rect 53880 115880 54120 115900
rect 54380 115880 54620 115900
rect 54880 115880 55120 115900
rect 55380 115880 55620 115900
rect 55880 115880 56120 115900
rect 56380 115880 56620 115900
rect 56880 115880 57120 115900
rect 57380 115880 57620 115900
rect 57880 115880 58000 115900
rect 14000 115620 14100 115880
rect 14400 115620 14600 115880
rect 14900 115620 15100 115880
rect 15400 115620 15600 115880
rect 15900 115620 16100 115880
rect 16400 115620 16600 115880
rect 16900 115620 17100 115880
rect 17400 115620 17600 115880
rect 17900 115620 18100 115880
rect 18400 115620 18600 115880
rect 18900 115620 19100 115880
rect 19400 115620 19600 115880
rect 19900 115620 20100 115880
rect 20400 115620 20600 115880
rect 20900 115620 21100 115880
rect 21400 115620 21600 115880
rect 21900 115620 22100 115880
rect 22400 115620 22600 115880
rect 22900 115620 23100 115880
rect 23400 115620 23600 115880
rect 23900 115620 24100 115880
rect 24400 115620 24600 115880
rect 24900 115620 25100 115880
rect 25400 115620 25600 115880
rect 25900 115620 26100 115880
rect 26400 115620 26600 115880
rect 26900 115620 27100 115880
rect 27400 115620 27600 115880
rect 27900 115620 28100 115880
rect 28400 115620 28600 115880
rect 28900 115620 29100 115880
rect 29400 115620 29600 115880
rect 29900 115620 30100 115880
rect 30400 115620 30600 115880
rect 30900 115620 31100 115880
rect 31400 115620 31600 115880
rect 31900 115620 32100 115880
rect 32400 115620 32600 115880
rect 32900 115620 33100 115880
rect 33400 115620 33600 115880
rect 33900 115620 34100 115880
rect 34400 115620 34600 115880
rect 34900 115620 35100 115880
rect 35400 115620 35600 115880
rect 35900 115620 36100 115880
rect 36400 115620 36600 115880
rect 36900 115620 37100 115880
rect 37400 115620 37600 115880
rect 37900 115620 38100 115880
rect 38400 115620 38600 115880
rect 38900 115620 39100 115880
rect 39400 115620 39600 115880
rect 39900 115620 40100 115880
rect 40400 115620 40600 115880
rect 40900 115620 41100 115880
rect 41400 115620 41600 115880
rect 41900 115620 42100 115880
rect 42400 115620 42600 115880
rect 42900 115620 43100 115880
rect 43400 115620 43600 115880
rect 43900 115620 44100 115880
rect 44400 115620 44600 115880
rect 44900 115620 45100 115880
rect 45400 115620 45600 115880
rect 45900 115620 46100 115880
rect 46400 115620 46600 115880
rect 46900 115620 47100 115880
rect 47400 115620 47600 115880
rect 47900 115620 48100 115880
rect 48400 115620 48600 115880
rect 48900 115620 49100 115880
rect 49400 115620 49600 115880
rect 49900 115620 50100 115880
rect 50400 115620 50600 115880
rect 50900 115620 51100 115880
rect 51400 115620 51600 115880
rect 51900 115620 52100 115880
rect 52400 115620 52600 115880
rect 52900 115620 53100 115880
rect 53400 115620 53600 115880
rect 53900 115620 54100 115880
rect 54400 115620 54600 115880
rect 54900 115620 55100 115880
rect 55400 115620 55600 115880
rect 55900 115620 56100 115880
rect 56400 115620 56600 115880
rect 56900 115620 57100 115880
rect 57400 115620 57600 115880
rect 57900 115620 58000 115880
rect 14000 115600 14120 115620
rect 14380 115600 14620 115620
rect 14880 115600 15120 115620
rect 15380 115600 15620 115620
rect 15880 115600 16120 115620
rect 16380 115600 16620 115620
rect 16880 115600 17120 115620
rect 17380 115600 17620 115620
rect 17880 115600 18120 115620
rect 18380 115600 18620 115620
rect 18880 115600 19120 115620
rect 19380 115600 19620 115620
rect 19880 115600 20120 115620
rect 20380 115600 20620 115620
rect 20880 115600 21120 115620
rect 21380 115600 21620 115620
rect 21880 115600 22120 115620
rect 22380 115600 22620 115620
rect 22880 115600 23120 115620
rect 23380 115600 23620 115620
rect 23880 115600 24120 115620
rect 24380 115600 24620 115620
rect 24880 115600 25120 115620
rect 25380 115600 25620 115620
rect 25880 115600 26120 115620
rect 26380 115600 26620 115620
rect 26880 115600 27120 115620
rect 27380 115600 27620 115620
rect 27880 115600 28120 115620
rect 28380 115600 28620 115620
rect 28880 115600 29120 115620
rect 29380 115600 29620 115620
rect 29880 115600 30120 115620
rect 30380 115600 30620 115620
rect 30880 115600 31120 115620
rect 31380 115600 31620 115620
rect 31880 115600 32120 115620
rect 32380 115600 32620 115620
rect 32880 115600 33120 115620
rect 33380 115600 33620 115620
rect 33880 115600 34120 115620
rect 34380 115600 34620 115620
rect 34880 115600 35120 115620
rect 35380 115600 35620 115620
rect 35880 115600 36120 115620
rect 36380 115600 36620 115620
rect 36880 115600 37120 115620
rect 37380 115600 37620 115620
rect 37880 115600 38120 115620
rect 38380 115600 38620 115620
rect 38880 115600 39120 115620
rect 39380 115600 39620 115620
rect 39880 115600 40120 115620
rect 40380 115600 40620 115620
rect 40880 115600 41120 115620
rect 41380 115600 41620 115620
rect 41880 115600 42120 115620
rect 42380 115600 42620 115620
rect 42880 115600 43120 115620
rect 43380 115600 43620 115620
rect 43880 115600 44120 115620
rect 44380 115600 44620 115620
rect 44880 115600 45120 115620
rect 45380 115600 45620 115620
rect 45880 115600 46120 115620
rect 46380 115600 46620 115620
rect 46880 115600 47120 115620
rect 47380 115600 47620 115620
rect 47880 115600 48120 115620
rect 48380 115600 48620 115620
rect 48880 115600 49120 115620
rect 49380 115600 49620 115620
rect 49880 115600 50120 115620
rect 50380 115600 50620 115620
rect 50880 115600 51120 115620
rect 51380 115600 51620 115620
rect 51880 115600 52120 115620
rect 52380 115600 52620 115620
rect 52880 115600 53120 115620
rect 53380 115600 53620 115620
rect 53880 115600 54120 115620
rect 54380 115600 54620 115620
rect 54880 115600 55120 115620
rect 55380 115600 55620 115620
rect 55880 115600 56120 115620
rect 56380 115600 56620 115620
rect 56880 115600 57120 115620
rect 57380 115600 57620 115620
rect 57880 115600 58000 115620
rect 14000 115400 58000 115600
rect 14000 115380 14120 115400
rect 14380 115380 14620 115400
rect 14880 115380 15120 115400
rect 15380 115380 15620 115400
rect 15880 115380 16120 115400
rect 16380 115380 16620 115400
rect 16880 115380 17120 115400
rect 17380 115380 17620 115400
rect 17880 115380 18120 115400
rect 18380 115380 18620 115400
rect 18880 115380 19120 115400
rect 19380 115380 19620 115400
rect 19880 115380 20120 115400
rect 20380 115380 20620 115400
rect 20880 115380 21120 115400
rect 21380 115380 21620 115400
rect 21880 115380 22120 115400
rect 22380 115380 22620 115400
rect 22880 115380 23120 115400
rect 23380 115380 23620 115400
rect 23880 115380 24120 115400
rect 24380 115380 24620 115400
rect 24880 115380 25120 115400
rect 25380 115380 25620 115400
rect 25880 115380 26120 115400
rect 26380 115380 26620 115400
rect 26880 115380 27120 115400
rect 27380 115380 27620 115400
rect 27880 115380 28120 115400
rect 28380 115380 28620 115400
rect 28880 115380 29120 115400
rect 29380 115380 29620 115400
rect 29880 115380 30120 115400
rect 30380 115380 30620 115400
rect 30880 115380 31120 115400
rect 31380 115380 31620 115400
rect 31880 115380 32120 115400
rect 32380 115380 32620 115400
rect 32880 115380 33120 115400
rect 33380 115380 33620 115400
rect 33880 115380 34120 115400
rect 34380 115380 34620 115400
rect 34880 115380 35120 115400
rect 35380 115380 35620 115400
rect 35880 115380 36120 115400
rect 36380 115380 36620 115400
rect 36880 115380 37120 115400
rect 37380 115380 37620 115400
rect 37880 115380 38120 115400
rect 38380 115380 38620 115400
rect 38880 115380 39120 115400
rect 39380 115380 39620 115400
rect 39880 115380 40120 115400
rect 40380 115380 40620 115400
rect 40880 115380 41120 115400
rect 41380 115380 41620 115400
rect 41880 115380 42120 115400
rect 42380 115380 42620 115400
rect 42880 115380 43120 115400
rect 43380 115380 43620 115400
rect 43880 115380 44120 115400
rect 44380 115380 44620 115400
rect 44880 115380 45120 115400
rect 45380 115380 45620 115400
rect 45880 115380 46120 115400
rect 46380 115380 46620 115400
rect 46880 115380 47120 115400
rect 47380 115380 47620 115400
rect 47880 115380 48120 115400
rect 48380 115380 48620 115400
rect 48880 115380 49120 115400
rect 49380 115380 49620 115400
rect 49880 115380 50120 115400
rect 50380 115380 50620 115400
rect 50880 115380 51120 115400
rect 51380 115380 51620 115400
rect 51880 115380 52120 115400
rect 52380 115380 52620 115400
rect 52880 115380 53120 115400
rect 53380 115380 53620 115400
rect 53880 115380 54120 115400
rect 54380 115380 54620 115400
rect 54880 115380 55120 115400
rect 55380 115380 55620 115400
rect 55880 115380 56120 115400
rect 56380 115380 56620 115400
rect 56880 115380 57120 115400
rect 57380 115380 57620 115400
rect 57880 115380 58000 115400
rect 14000 115120 14100 115380
rect 14400 115120 14600 115380
rect 14900 115120 15100 115380
rect 15400 115120 15600 115380
rect 15900 115120 16100 115380
rect 16400 115120 16600 115380
rect 16900 115120 17100 115380
rect 17400 115120 17600 115380
rect 17900 115120 18100 115380
rect 18400 115120 18600 115380
rect 18900 115120 19100 115380
rect 19400 115120 19600 115380
rect 19900 115120 20100 115380
rect 20400 115120 20600 115380
rect 20900 115120 21100 115380
rect 21400 115120 21600 115380
rect 21900 115120 22100 115380
rect 22400 115120 22600 115380
rect 22900 115120 23100 115380
rect 23400 115120 23600 115380
rect 23900 115120 24100 115380
rect 24400 115120 24600 115380
rect 24900 115120 25100 115380
rect 25400 115120 25600 115380
rect 25900 115120 26100 115380
rect 26400 115120 26600 115380
rect 26900 115120 27100 115380
rect 27400 115120 27600 115380
rect 27900 115120 28100 115380
rect 28400 115120 28600 115380
rect 28900 115120 29100 115380
rect 29400 115120 29600 115380
rect 29900 115120 30100 115380
rect 30400 115120 30600 115380
rect 30900 115120 31100 115380
rect 31400 115120 31600 115380
rect 31900 115120 32100 115380
rect 32400 115120 32600 115380
rect 32900 115120 33100 115380
rect 33400 115120 33600 115380
rect 33900 115120 34100 115380
rect 34400 115120 34600 115380
rect 34900 115120 35100 115380
rect 35400 115120 35600 115380
rect 35900 115120 36100 115380
rect 36400 115120 36600 115380
rect 36900 115120 37100 115380
rect 37400 115120 37600 115380
rect 37900 115120 38100 115380
rect 38400 115120 38600 115380
rect 38900 115120 39100 115380
rect 39400 115120 39600 115380
rect 39900 115120 40100 115380
rect 40400 115120 40600 115380
rect 40900 115120 41100 115380
rect 41400 115120 41600 115380
rect 41900 115120 42100 115380
rect 42400 115120 42600 115380
rect 42900 115120 43100 115380
rect 43400 115120 43600 115380
rect 43900 115120 44100 115380
rect 44400 115120 44600 115380
rect 44900 115120 45100 115380
rect 45400 115120 45600 115380
rect 45900 115120 46100 115380
rect 46400 115120 46600 115380
rect 46900 115120 47100 115380
rect 47400 115120 47600 115380
rect 47900 115120 48100 115380
rect 48400 115120 48600 115380
rect 48900 115120 49100 115380
rect 49400 115120 49600 115380
rect 49900 115120 50100 115380
rect 50400 115120 50600 115380
rect 50900 115120 51100 115380
rect 51400 115120 51600 115380
rect 51900 115120 52100 115380
rect 52400 115120 52600 115380
rect 52900 115120 53100 115380
rect 53400 115120 53600 115380
rect 53900 115120 54100 115380
rect 54400 115120 54600 115380
rect 54900 115120 55100 115380
rect 55400 115120 55600 115380
rect 55900 115120 56100 115380
rect 56400 115120 56600 115380
rect 56900 115120 57100 115380
rect 57400 115120 57600 115380
rect 57900 115120 58000 115380
rect 14000 115100 14120 115120
rect 14380 115100 14620 115120
rect 14880 115100 15120 115120
rect 15380 115100 15620 115120
rect 15880 115100 16120 115120
rect 16380 115100 16620 115120
rect 16880 115100 17120 115120
rect 17380 115100 17620 115120
rect 17880 115100 18120 115120
rect 18380 115100 18620 115120
rect 18880 115100 19120 115120
rect 19380 115100 19620 115120
rect 19880 115100 20120 115120
rect 20380 115100 20620 115120
rect 20880 115100 21120 115120
rect 21380 115100 21620 115120
rect 21880 115100 22120 115120
rect 22380 115100 22620 115120
rect 22880 115100 23120 115120
rect 23380 115100 23620 115120
rect 23880 115100 24120 115120
rect 24380 115100 24620 115120
rect 24880 115100 25120 115120
rect 25380 115100 25620 115120
rect 25880 115100 26120 115120
rect 26380 115100 26620 115120
rect 26880 115100 27120 115120
rect 27380 115100 27620 115120
rect 27880 115100 28120 115120
rect 28380 115100 28620 115120
rect 28880 115100 29120 115120
rect 29380 115100 29620 115120
rect 29880 115100 30120 115120
rect 30380 115100 30620 115120
rect 30880 115100 31120 115120
rect 31380 115100 31620 115120
rect 31880 115100 32120 115120
rect 32380 115100 32620 115120
rect 32880 115100 33120 115120
rect 33380 115100 33620 115120
rect 33880 115100 34120 115120
rect 34380 115100 34620 115120
rect 34880 115100 35120 115120
rect 35380 115100 35620 115120
rect 35880 115100 36120 115120
rect 36380 115100 36620 115120
rect 36880 115100 37120 115120
rect 37380 115100 37620 115120
rect 37880 115100 38120 115120
rect 38380 115100 38620 115120
rect 38880 115100 39120 115120
rect 39380 115100 39620 115120
rect 39880 115100 40120 115120
rect 40380 115100 40620 115120
rect 40880 115100 41120 115120
rect 41380 115100 41620 115120
rect 41880 115100 42120 115120
rect 42380 115100 42620 115120
rect 42880 115100 43120 115120
rect 43380 115100 43620 115120
rect 43880 115100 44120 115120
rect 44380 115100 44620 115120
rect 44880 115100 45120 115120
rect 45380 115100 45620 115120
rect 45880 115100 46120 115120
rect 46380 115100 46620 115120
rect 46880 115100 47120 115120
rect 47380 115100 47620 115120
rect 47880 115100 48120 115120
rect 48380 115100 48620 115120
rect 48880 115100 49120 115120
rect 49380 115100 49620 115120
rect 49880 115100 50120 115120
rect 50380 115100 50620 115120
rect 50880 115100 51120 115120
rect 51380 115100 51620 115120
rect 51880 115100 52120 115120
rect 52380 115100 52620 115120
rect 52880 115100 53120 115120
rect 53380 115100 53620 115120
rect 53880 115100 54120 115120
rect 54380 115100 54620 115120
rect 54880 115100 55120 115120
rect 55380 115100 55620 115120
rect 55880 115100 56120 115120
rect 56380 115100 56620 115120
rect 56880 115100 57120 115120
rect 57380 115100 57620 115120
rect 57880 115100 58000 115120
rect 14000 114900 58000 115100
rect 14000 114880 14120 114900
rect 14380 114880 14620 114900
rect 14880 114880 15120 114900
rect 15380 114880 15620 114900
rect 15880 114880 16120 114900
rect 16380 114880 16620 114900
rect 16880 114880 17120 114900
rect 17380 114880 17620 114900
rect 17880 114880 18120 114900
rect 18380 114880 18620 114900
rect 18880 114880 19120 114900
rect 19380 114880 19620 114900
rect 19880 114880 20120 114900
rect 20380 114880 20620 114900
rect 20880 114880 21120 114900
rect 21380 114880 21620 114900
rect 21880 114880 22120 114900
rect 22380 114880 22620 114900
rect 22880 114880 23120 114900
rect 23380 114880 23620 114900
rect 23880 114880 24120 114900
rect 24380 114880 24620 114900
rect 24880 114880 25120 114900
rect 25380 114880 25620 114900
rect 25880 114880 26120 114900
rect 26380 114880 26620 114900
rect 26880 114880 27120 114900
rect 27380 114880 27620 114900
rect 27880 114880 28120 114900
rect 28380 114880 28620 114900
rect 28880 114880 29120 114900
rect 29380 114880 29620 114900
rect 29880 114880 30120 114900
rect 30380 114880 30620 114900
rect 30880 114880 31120 114900
rect 31380 114880 31620 114900
rect 31880 114880 32120 114900
rect 32380 114880 32620 114900
rect 32880 114880 33120 114900
rect 33380 114880 33620 114900
rect 33880 114880 34120 114900
rect 34380 114880 34620 114900
rect 34880 114880 35120 114900
rect 35380 114880 35620 114900
rect 35880 114880 36120 114900
rect 36380 114880 36620 114900
rect 36880 114880 37120 114900
rect 37380 114880 37620 114900
rect 37880 114880 38120 114900
rect 38380 114880 38620 114900
rect 38880 114880 39120 114900
rect 39380 114880 39620 114900
rect 39880 114880 40120 114900
rect 40380 114880 40620 114900
rect 40880 114880 41120 114900
rect 41380 114880 41620 114900
rect 41880 114880 42120 114900
rect 42380 114880 42620 114900
rect 42880 114880 43120 114900
rect 43380 114880 43620 114900
rect 43880 114880 44120 114900
rect 44380 114880 44620 114900
rect 44880 114880 45120 114900
rect 45380 114880 45620 114900
rect 45880 114880 46120 114900
rect 46380 114880 46620 114900
rect 46880 114880 47120 114900
rect 47380 114880 47620 114900
rect 47880 114880 48120 114900
rect 48380 114880 48620 114900
rect 48880 114880 49120 114900
rect 49380 114880 49620 114900
rect 49880 114880 50120 114900
rect 50380 114880 50620 114900
rect 50880 114880 51120 114900
rect 51380 114880 51620 114900
rect 51880 114880 52120 114900
rect 52380 114880 52620 114900
rect 52880 114880 53120 114900
rect 53380 114880 53620 114900
rect 53880 114880 54120 114900
rect 54380 114880 54620 114900
rect 54880 114880 55120 114900
rect 55380 114880 55620 114900
rect 55880 114880 56120 114900
rect 56380 114880 56620 114900
rect 56880 114880 57120 114900
rect 57380 114880 57620 114900
rect 57880 114880 58000 114900
rect 14000 114620 14100 114880
rect 14400 114620 14600 114880
rect 14900 114620 15100 114880
rect 15400 114620 15600 114880
rect 15900 114620 16100 114880
rect 16400 114620 16600 114880
rect 16900 114620 17100 114880
rect 17400 114620 17600 114880
rect 17900 114620 18100 114880
rect 18400 114620 18600 114880
rect 18900 114620 19100 114880
rect 19400 114620 19600 114880
rect 19900 114620 20100 114880
rect 20400 114620 20600 114880
rect 20900 114620 21100 114880
rect 21400 114620 21600 114880
rect 21900 114620 22100 114880
rect 22400 114620 22600 114880
rect 22900 114620 23100 114880
rect 23400 114620 23600 114880
rect 23900 114620 24100 114880
rect 24400 114620 24600 114880
rect 24900 114620 25100 114880
rect 25400 114620 25600 114880
rect 25900 114620 26100 114880
rect 26400 114620 26600 114880
rect 26900 114620 27100 114880
rect 27400 114620 27600 114880
rect 27900 114620 28100 114880
rect 28400 114620 28600 114880
rect 28900 114620 29100 114880
rect 29400 114620 29600 114880
rect 29900 114620 30100 114880
rect 30400 114620 30600 114880
rect 30900 114620 31100 114880
rect 31400 114620 31600 114880
rect 31900 114620 32100 114880
rect 32400 114620 32600 114880
rect 32900 114620 33100 114880
rect 33400 114620 33600 114880
rect 33900 114620 34100 114880
rect 34400 114620 34600 114880
rect 34900 114620 35100 114880
rect 35400 114620 35600 114880
rect 35900 114620 36100 114880
rect 36400 114620 36600 114880
rect 36900 114620 37100 114880
rect 37400 114620 37600 114880
rect 37900 114620 38100 114880
rect 38400 114620 38600 114880
rect 38900 114620 39100 114880
rect 39400 114620 39600 114880
rect 39900 114620 40100 114880
rect 40400 114620 40600 114880
rect 40900 114620 41100 114880
rect 41400 114620 41600 114880
rect 41900 114620 42100 114880
rect 42400 114620 42600 114880
rect 42900 114620 43100 114880
rect 43400 114620 43600 114880
rect 43900 114620 44100 114880
rect 44400 114620 44600 114880
rect 44900 114620 45100 114880
rect 45400 114620 45600 114880
rect 45900 114620 46100 114880
rect 46400 114620 46600 114880
rect 46900 114620 47100 114880
rect 47400 114620 47600 114880
rect 47900 114620 48100 114880
rect 48400 114620 48600 114880
rect 48900 114620 49100 114880
rect 49400 114620 49600 114880
rect 49900 114620 50100 114880
rect 50400 114620 50600 114880
rect 50900 114620 51100 114880
rect 51400 114620 51600 114880
rect 51900 114620 52100 114880
rect 52400 114620 52600 114880
rect 52900 114620 53100 114880
rect 53400 114620 53600 114880
rect 53900 114620 54100 114880
rect 54400 114620 54600 114880
rect 54900 114620 55100 114880
rect 55400 114620 55600 114880
rect 55900 114620 56100 114880
rect 56400 114620 56600 114880
rect 56900 114620 57100 114880
rect 57400 114620 57600 114880
rect 57900 114620 58000 114880
rect 14000 114600 14120 114620
rect 14380 114600 14620 114620
rect 14880 114600 15120 114620
rect 15380 114600 15620 114620
rect 15880 114600 16120 114620
rect 16380 114600 16620 114620
rect 16880 114600 17120 114620
rect 17380 114600 17620 114620
rect 17880 114600 18120 114620
rect 18380 114600 18620 114620
rect 18880 114600 19120 114620
rect 19380 114600 19620 114620
rect 19880 114600 20120 114620
rect 20380 114600 20620 114620
rect 20880 114600 21120 114620
rect 21380 114600 21620 114620
rect 21880 114600 22120 114620
rect 22380 114600 22620 114620
rect 22880 114600 23120 114620
rect 23380 114600 23620 114620
rect 23880 114600 24120 114620
rect 24380 114600 24620 114620
rect 24880 114600 25120 114620
rect 25380 114600 25620 114620
rect 25880 114600 26120 114620
rect 26380 114600 26620 114620
rect 26880 114600 27120 114620
rect 27380 114600 27620 114620
rect 27880 114600 28120 114620
rect 28380 114600 28620 114620
rect 28880 114600 29120 114620
rect 29380 114600 29620 114620
rect 29880 114600 30120 114620
rect 30380 114600 30620 114620
rect 30880 114600 31120 114620
rect 31380 114600 31620 114620
rect 31880 114600 32120 114620
rect 32380 114600 32620 114620
rect 32880 114600 33120 114620
rect 33380 114600 33620 114620
rect 33880 114600 34120 114620
rect 34380 114600 34620 114620
rect 34880 114600 35120 114620
rect 35380 114600 35620 114620
rect 35880 114600 36120 114620
rect 36380 114600 36620 114620
rect 36880 114600 37120 114620
rect 37380 114600 37620 114620
rect 37880 114600 38120 114620
rect 38380 114600 38620 114620
rect 38880 114600 39120 114620
rect 39380 114600 39620 114620
rect 39880 114600 40120 114620
rect 40380 114600 40620 114620
rect 40880 114600 41120 114620
rect 41380 114600 41620 114620
rect 41880 114600 42120 114620
rect 42380 114600 42620 114620
rect 42880 114600 43120 114620
rect 43380 114600 43620 114620
rect 43880 114600 44120 114620
rect 44380 114600 44620 114620
rect 44880 114600 45120 114620
rect 45380 114600 45620 114620
rect 45880 114600 46120 114620
rect 46380 114600 46620 114620
rect 46880 114600 47120 114620
rect 47380 114600 47620 114620
rect 47880 114600 48120 114620
rect 48380 114600 48620 114620
rect 48880 114600 49120 114620
rect 49380 114600 49620 114620
rect 49880 114600 50120 114620
rect 50380 114600 50620 114620
rect 50880 114600 51120 114620
rect 51380 114600 51620 114620
rect 51880 114600 52120 114620
rect 52380 114600 52620 114620
rect 52880 114600 53120 114620
rect 53380 114600 53620 114620
rect 53880 114600 54120 114620
rect 54380 114600 54620 114620
rect 54880 114600 55120 114620
rect 55380 114600 55620 114620
rect 55880 114600 56120 114620
rect 56380 114600 56620 114620
rect 56880 114600 57120 114620
rect 57380 114600 57620 114620
rect 57880 114600 58000 114620
rect 14000 114400 58000 114600
rect 14000 114380 14120 114400
rect 14380 114380 14620 114400
rect 14880 114380 15120 114400
rect 15380 114380 15620 114400
rect 15880 114380 16120 114400
rect 16380 114380 16620 114400
rect 16880 114380 17120 114400
rect 17380 114380 17620 114400
rect 17880 114380 18120 114400
rect 18380 114380 18620 114400
rect 18880 114380 19120 114400
rect 19380 114380 19620 114400
rect 19880 114380 20120 114400
rect 20380 114380 20620 114400
rect 20880 114380 21120 114400
rect 21380 114380 21620 114400
rect 21880 114380 22120 114400
rect 22380 114380 22620 114400
rect 22880 114380 23120 114400
rect 23380 114380 23620 114400
rect 23880 114380 24120 114400
rect 24380 114380 24620 114400
rect 24880 114380 25120 114400
rect 25380 114380 25620 114400
rect 25880 114380 26120 114400
rect 26380 114380 26620 114400
rect 26880 114380 27120 114400
rect 27380 114380 27620 114400
rect 27880 114380 28120 114400
rect 28380 114380 28620 114400
rect 28880 114380 29120 114400
rect 29380 114380 29620 114400
rect 29880 114380 30120 114400
rect 30380 114380 30620 114400
rect 30880 114380 31120 114400
rect 31380 114380 31620 114400
rect 31880 114380 32120 114400
rect 32380 114380 32620 114400
rect 32880 114380 33120 114400
rect 33380 114380 33620 114400
rect 33880 114380 34120 114400
rect 34380 114380 34620 114400
rect 34880 114380 35120 114400
rect 35380 114380 35620 114400
rect 35880 114380 36120 114400
rect 36380 114380 36620 114400
rect 36880 114380 37120 114400
rect 37380 114380 37620 114400
rect 37880 114380 38120 114400
rect 38380 114380 38620 114400
rect 38880 114380 39120 114400
rect 39380 114380 39620 114400
rect 39880 114380 40120 114400
rect 40380 114380 40620 114400
rect 40880 114380 41120 114400
rect 41380 114380 41620 114400
rect 41880 114380 42120 114400
rect 42380 114380 42620 114400
rect 42880 114380 43120 114400
rect 43380 114380 43620 114400
rect 43880 114380 44120 114400
rect 44380 114380 44620 114400
rect 44880 114380 45120 114400
rect 45380 114380 45620 114400
rect 45880 114380 46120 114400
rect 46380 114380 46620 114400
rect 46880 114380 47120 114400
rect 47380 114380 47620 114400
rect 47880 114380 48120 114400
rect 48380 114380 48620 114400
rect 48880 114380 49120 114400
rect 49380 114380 49620 114400
rect 49880 114380 50120 114400
rect 50380 114380 50620 114400
rect 50880 114380 51120 114400
rect 51380 114380 51620 114400
rect 51880 114380 52120 114400
rect 52380 114380 52620 114400
rect 52880 114380 53120 114400
rect 53380 114380 53620 114400
rect 53880 114380 54120 114400
rect 54380 114380 54620 114400
rect 54880 114380 55120 114400
rect 55380 114380 55620 114400
rect 55880 114380 56120 114400
rect 56380 114380 56620 114400
rect 56880 114380 57120 114400
rect 57380 114380 57620 114400
rect 57880 114380 58000 114400
rect 14000 114120 14100 114380
rect 14400 114120 14600 114380
rect 14900 114120 15100 114380
rect 15400 114120 15600 114380
rect 15900 114120 16100 114380
rect 16400 114120 16600 114380
rect 16900 114120 17100 114380
rect 17400 114120 17600 114380
rect 17900 114120 18100 114380
rect 18400 114120 18600 114380
rect 18900 114120 19100 114380
rect 19400 114120 19600 114380
rect 19900 114120 20100 114380
rect 20400 114120 20600 114380
rect 20900 114120 21100 114380
rect 21400 114120 21600 114380
rect 21900 114120 22100 114380
rect 22400 114120 22600 114380
rect 22900 114120 23100 114380
rect 23400 114120 23600 114380
rect 23900 114120 24100 114380
rect 24400 114120 24600 114380
rect 24900 114120 25100 114380
rect 25400 114120 25600 114380
rect 25900 114120 26100 114380
rect 26400 114120 26600 114380
rect 26900 114120 27100 114380
rect 27400 114120 27600 114380
rect 27900 114120 28100 114380
rect 28400 114120 28600 114380
rect 28900 114120 29100 114380
rect 29400 114120 29600 114380
rect 29900 114120 30100 114380
rect 30400 114120 30600 114380
rect 30900 114120 31100 114380
rect 31400 114120 31600 114380
rect 31900 114120 32100 114380
rect 32400 114120 32600 114380
rect 32900 114120 33100 114380
rect 33400 114120 33600 114380
rect 33900 114120 34100 114380
rect 34400 114120 34600 114380
rect 34900 114120 35100 114380
rect 35400 114120 35600 114380
rect 35900 114120 36100 114380
rect 36400 114120 36600 114380
rect 36900 114120 37100 114380
rect 37400 114120 37600 114380
rect 37900 114120 38100 114380
rect 38400 114120 38600 114380
rect 38900 114120 39100 114380
rect 39400 114120 39600 114380
rect 39900 114120 40100 114380
rect 40400 114120 40600 114380
rect 40900 114120 41100 114380
rect 41400 114120 41600 114380
rect 41900 114120 42100 114380
rect 42400 114120 42600 114380
rect 42900 114120 43100 114380
rect 43400 114120 43600 114380
rect 43900 114120 44100 114380
rect 44400 114120 44600 114380
rect 44900 114120 45100 114380
rect 45400 114120 45600 114380
rect 45900 114120 46100 114380
rect 46400 114120 46600 114380
rect 46900 114120 47100 114380
rect 47400 114120 47600 114380
rect 47900 114120 48100 114380
rect 48400 114120 48600 114380
rect 48900 114120 49100 114380
rect 49400 114120 49600 114380
rect 49900 114120 50100 114380
rect 50400 114120 50600 114380
rect 50900 114120 51100 114380
rect 51400 114120 51600 114380
rect 51900 114120 52100 114380
rect 52400 114120 52600 114380
rect 52900 114120 53100 114380
rect 53400 114120 53600 114380
rect 53900 114120 54100 114380
rect 54400 114120 54600 114380
rect 54900 114120 55100 114380
rect 55400 114120 55600 114380
rect 55900 114120 56100 114380
rect 56400 114120 56600 114380
rect 56900 114120 57100 114380
rect 57400 114120 57600 114380
rect 57900 114120 58000 114380
rect 14000 114100 14120 114120
rect 14380 114100 14620 114120
rect 14880 114100 15120 114120
rect 15380 114100 15620 114120
rect 15880 114100 16120 114120
rect 16380 114100 16620 114120
rect 16880 114100 17120 114120
rect 17380 114100 17620 114120
rect 17880 114100 18120 114120
rect 18380 114100 18620 114120
rect 18880 114100 19120 114120
rect 19380 114100 19620 114120
rect 19880 114100 20120 114120
rect 20380 114100 20620 114120
rect 20880 114100 21120 114120
rect 21380 114100 21620 114120
rect 21880 114100 22120 114120
rect 22380 114100 22620 114120
rect 22880 114100 23120 114120
rect 23380 114100 23620 114120
rect 23880 114100 24120 114120
rect 24380 114100 24620 114120
rect 24880 114100 25120 114120
rect 25380 114100 25620 114120
rect 25880 114100 26120 114120
rect 26380 114100 26620 114120
rect 26880 114100 27120 114120
rect 27380 114100 27620 114120
rect 27880 114100 28120 114120
rect 28380 114100 28620 114120
rect 28880 114100 29120 114120
rect 29380 114100 29620 114120
rect 29880 114100 30120 114120
rect 30380 114100 30620 114120
rect 30880 114100 31120 114120
rect 31380 114100 31620 114120
rect 31880 114100 32120 114120
rect 32380 114100 32620 114120
rect 32880 114100 33120 114120
rect 33380 114100 33620 114120
rect 33880 114100 34120 114120
rect 34380 114100 34620 114120
rect 34880 114100 35120 114120
rect 35380 114100 35620 114120
rect 35880 114100 36120 114120
rect 36380 114100 36620 114120
rect 36880 114100 37120 114120
rect 37380 114100 37620 114120
rect 37880 114100 38120 114120
rect 38380 114100 38620 114120
rect 38880 114100 39120 114120
rect 39380 114100 39620 114120
rect 39880 114100 40120 114120
rect 40380 114100 40620 114120
rect 40880 114100 41120 114120
rect 41380 114100 41620 114120
rect 41880 114100 42120 114120
rect 42380 114100 42620 114120
rect 42880 114100 43120 114120
rect 43380 114100 43620 114120
rect 43880 114100 44120 114120
rect 44380 114100 44620 114120
rect 44880 114100 45120 114120
rect 45380 114100 45620 114120
rect 45880 114100 46120 114120
rect 46380 114100 46620 114120
rect 46880 114100 47120 114120
rect 47380 114100 47620 114120
rect 47880 114100 48120 114120
rect 48380 114100 48620 114120
rect 48880 114100 49120 114120
rect 49380 114100 49620 114120
rect 49880 114100 50120 114120
rect 50380 114100 50620 114120
rect 50880 114100 51120 114120
rect 51380 114100 51620 114120
rect 51880 114100 52120 114120
rect 52380 114100 52620 114120
rect 52880 114100 53120 114120
rect 53380 114100 53620 114120
rect 53880 114100 54120 114120
rect 54380 114100 54620 114120
rect 54880 114100 55120 114120
rect 55380 114100 55620 114120
rect 55880 114100 56120 114120
rect 56380 114100 56620 114120
rect 56880 114100 57120 114120
rect 57380 114100 57620 114120
rect 57880 114100 58000 114120
rect 14000 114000 58000 114100
rect 118000 121900 142000 122000
rect 118000 121880 118120 121900
rect 118380 121880 118620 121900
rect 118880 121880 119120 121900
rect 119380 121880 119620 121900
rect 119880 121880 120120 121900
rect 120380 121880 120620 121900
rect 120880 121880 121120 121900
rect 121380 121880 121620 121900
rect 121880 121880 122120 121900
rect 122380 121880 122620 121900
rect 122880 121880 123120 121900
rect 123380 121880 123620 121900
rect 123880 121880 124120 121900
rect 124380 121880 124620 121900
rect 124880 121880 125120 121900
rect 125380 121880 125620 121900
rect 125880 121880 126120 121900
rect 126380 121880 126620 121900
rect 126880 121880 127120 121900
rect 127380 121880 127620 121900
rect 127880 121880 128120 121900
rect 128380 121880 128620 121900
rect 128880 121880 129120 121900
rect 129380 121880 129620 121900
rect 129880 121880 130120 121900
rect 130380 121880 130620 121900
rect 130880 121880 131120 121900
rect 131380 121880 131620 121900
rect 131880 121880 132120 121900
rect 132380 121880 132620 121900
rect 132880 121880 133120 121900
rect 133380 121880 133620 121900
rect 133880 121880 134120 121900
rect 134380 121880 134620 121900
rect 134880 121880 135120 121900
rect 135380 121880 135620 121900
rect 135880 121880 136120 121900
rect 136380 121880 136620 121900
rect 136880 121880 137120 121900
rect 137380 121880 137620 121900
rect 137880 121880 138120 121900
rect 138380 121880 138620 121900
rect 138880 121880 139120 121900
rect 139380 121880 139620 121900
rect 139880 121880 140120 121900
rect 140380 121880 140620 121900
rect 140880 121880 141120 121900
rect 141380 121880 141620 121900
rect 141880 121880 142000 121900
rect 118000 121620 118100 121880
rect 118400 121620 118600 121880
rect 118900 121620 119100 121880
rect 119400 121620 119600 121880
rect 119900 121620 120100 121880
rect 120400 121620 120600 121880
rect 120900 121620 121100 121880
rect 121400 121620 121600 121880
rect 121900 121620 122100 121880
rect 122400 121620 122600 121880
rect 122900 121620 123100 121880
rect 123400 121620 123600 121880
rect 123900 121620 124100 121880
rect 124400 121620 124600 121880
rect 124900 121620 125100 121880
rect 125400 121620 125600 121880
rect 125900 121620 126100 121880
rect 126400 121620 126600 121880
rect 126900 121620 127100 121880
rect 127400 121620 127600 121880
rect 127900 121620 128100 121880
rect 128400 121620 128600 121880
rect 128900 121620 129100 121880
rect 129400 121620 129600 121880
rect 129900 121620 130100 121880
rect 130400 121620 130600 121880
rect 130900 121620 131100 121880
rect 131400 121620 131600 121880
rect 131900 121620 132100 121880
rect 132400 121620 132600 121880
rect 132900 121620 133100 121880
rect 133400 121620 133600 121880
rect 133900 121620 134100 121880
rect 134400 121620 134600 121880
rect 134900 121620 135100 121880
rect 135400 121620 135600 121880
rect 135900 121620 136100 121880
rect 136400 121620 136600 121880
rect 136900 121620 137100 121880
rect 137400 121620 137600 121880
rect 137900 121620 138100 121880
rect 138400 121620 138600 121880
rect 138900 121620 139100 121880
rect 139400 121620 139600 121880
rect 139900 121620 140100 121880
rect 140400 121620 140600 121880
rect 140900 121620 141100 121880
rect 141400 121620 141600 121880
rect 141900 121620 142000 121880
rect 118000 121600 118120 121620
rect 118380 121600 118620 121620
rect 118880 121600 119120 121620
rect 119380 121600 119620 121620
rect 119880 121600 120120 121620
rect 120380 121600 120620 121620
rect 120880 121600 121120 121620
rect 121380 121600 121620 121620
rect 121880 121600 122120 121620
rect 122380 121600 122620 121620
rect 122880 121600 123120 121620
rect 123380 121600 123620 121620
rect 123880 121600 124120 121620
rect 124380 121600 124620 121620
rect 124880 121600 125120 121620
rect 125380 121600 125620 121620
rect 125880 121600 126120 121620
rect 126380 121600 126620 121620
rect 126880 121600 127120 121620
rect 127380 121600 127620 121620
rect 127880 121600 128120 121620
rect 128380 121600 128620 121620
rect 128880 121600 129120 121620
rect 129380 121600 129620 121620
rect 129880 121600 130120 121620
rect 130380 121600 130620 121620
rect 130880 121600 131120 121620
rect 131380 121600 131620 121620
rect 131880 121600 132120 121620
rect 132380 121600 132620 121620
rect 132880 121600 133120 121620
rect 133380 121600 133620 121620
rect 133880 121600 134120 121620
rect 134380 121600 134620 121620
rect 134880 121600 135120 121620
rect 135380 121600 135620 121620
rect 135880 121600 136120 121620
rect 136380 121600 136620 121620
rect 136880 121600 137120 121620
rect 137380 121600 137620 121620
rect 137880 121600 138120 121620
rect 138380 121600 138620 121620
rect 138880 121600 139120 121620
rect 139380 121600 139620 121620
rect 139880 121600 140120 121620
rect 140380 121600 140620 121620
rect 140880 121600 141120 121620
rect 141380 121600 141620 121620
rect 141880 121600 142000 121620
rect 118000 121400 142000 121600
rect 118000 121380 118120 121400
rect 118380 121380 118620 121400
rect 118880 121380 119120 121400
rect 119380 121380 119620 121400
rect 119880 121380 120120 121400
rect 120380 121380 120620 121400
rect 120880 121380 121120 121400
rect 121380 121380 121620 121400
rect 121880 121380 122120 121400
rect 122380 121380 122620 121400
rect 122880 121380 123120 121400
rect 123380 121380 123620 121400
rect 123880 121380 124120 121400
rect 124380 121380 124620 121400
rect 124880 121380 125120 121400
rect 125380 121380 125620 121400
rect 125880 121380 126120 121400
rect 126380 121380 126620 121400
rect 126880 121380 127120 121400
rect 127380 121380 127620 121400
rect 127880 121380 128120 121400
rect 128380 121380 128620 121400
rect 128880 121380 129120 121400
rect 129380 121380 129620 121400
rect 129880 121380 130120 121400
rect 130380 121380 130620 121400
rect 130880 121380 131120 121400
rect 131380 121380 131620 121400
rect 131880 121380 132120 121400
rect 132380 121380 132620 121400
rect 132880 121380 133120 121400
rect 133380 121380 133620 121400
rect 133880 121380 134120 121400
rect 134380 121380 134620 121400
rect 134880 121380 135120 121400
rect 135380 121380 135620 121400
rect 135880 121380 136120 121400
rect 136380 121380 136620 121400
rect 136880 121380 137120 121400
rect 137380 121380 137620 121400
rect 137880 121380 138120 121400
rect 138380 121380 138620 121400
rect 138880 121380 139120 121400
rect 139380 121380 139620 121400
rect 139880 121380 140120 121400
rect 140380 121380 140620 121400
rect 140880 121380 141120 121400
rect 141380 121380 141620 121400
rect 141880 121380 142000 121400
rect 118000 121120 118100 121380
rect 118400 121120 118600 121380
rect 118900 121120 119100 121380
rect 119400 121120 119600 121380
rect 119900 121120 120100 121380
rect 120400 121120 120600 121380
rect 120900 121120 121100 121380
rect 121400 121120 121600 121380
rect 121900 121120 122100 121380
rect 122400 121120 122600 121380
rect 122900 121120 123100 121380
rect 123400 121120 123600 121380
rect 123900 121120 124100 121380
rect 124400 121120 124600 121380
rect 124900 121120 125100 121380
rect 125400 121120 125600 121380
rect 125900 121120 126100 121380
rect 126400 121120 126600 121380
rect 126900 121120 127100 121380
rect 127400 121120 127600 121380
rect 127900 121120 128100 121380
rect 128400 121120 128600 121380
rect 128900 121120 129100 121380
rect 129400 121120 129600 121380
rect 129900 121120 130100 121380
rect 130400 121120 130600 121380
rect 130900 121120 131100 121380
rect 131400 121120 131600 121380
rect 131900 121120 132100 121380
rect 132400 121120 132600 121380
rect 132900 121120 133100 121380
rect 133400 121120 133600 121380
rect 133900 121120 134100 121380
rect 134400 121120 134600 121380
rect 134900 121120 135100 121380
rect 135400 121120 135600 121380
rect 135900 121120 136100 121380
rect 136400 121120 136600 121380
rect 136900 121120 137100 121380
rect 137400 121120 137600 121380
rect 137900 121120 138100 121380
rect 138400 121120 138600 121380
rect 138900 121120 139100 121380
rect 139400 121120 139600 121380
rect 139900 121120 140100 121380
rect 140400 121120 140600 121380
rect 140900 121120 141100 121380
rect 141400 121120 141600 121380
rect 141900 121120 142000 121380
rect 118000 121100 118120 121120
rect 118380 121100 118620 121120
rect 118880 121100 119120 121120
rect 119380 121100 119620 121120
rect 119880 121100 120120 121120
rect 120380 121100 120620 121120
rect 120880 121100 121120 121120
rect 121380 121100 121620 121120
rect 121880 121100 122120 121120
rect 122380 121100 122620 121120
rect 122880 121100 123120 121120
rect 123380 121100 123620 121120
rect 123880 121100 124120 121120
rect 124380 121100 124620 121120
rect 124880 121100 125120 121120
rect 125380 121100 125620 121120
rect 125880 121100 126120 121120
rect 126380 121100 126620 121120
rect 126880 121100 127120 121120
rect 127380 121100 127620 121120
rect 127880 121100 128120 121120
rect 128380 121100 128620 121120
rect 128880 121100 129120 121120
rect 129380 121100 129620 121120
rect 129880 121100 130120 121120
rect 130380 121100 130620 121120
rect 130880 121100 131120 121120
rect 131380 121100 131620 121120
rect 131880 121100 132120 121120
rect 132380 121100 132620 121120
rect 132880 121100 133120 121120
rect 133380 121100 133620 121120
rect 133880 121100 134120 121120
rect 134380 121100 134620 121120
rect 134880 121100 135120 121120
rect 135380 121100 135620 121120
rect 135880 121100 136120 121120
rect 136380 121100 136620 121120
rect 136880 121100 137120 121120
rect 137380 121100 137620 121120
rect 137880 121100 138120 121120
rect 138380 121100 138620 121120
rect 138880 121100 139120 121120
rect 139380 121100 139620 121120
rect 139880 121100 140120 121120
rect 140380 121100 140620 121120
rect 140880 121100 141120 121120
rect 141380 121100 141620 121120
rect 141880 121100 142000 121120
rect 118000 120900 142000 121100
rect 118000 120880 118120 120900
rect 118380 120880 118620 120900
rect 118880 120880 119120 120900
rect 119380 120880 119620 120900
rect 119880 120880 120120 120900
rect 120380 120880 120620 120900
rect 120880 120880 121120 120900
rect 121380 120880 121620 120900
rect 121880 120880 122120 120900
rect 122380 120880 122620 120900
rect 122880 120880 123120 120900
rect 123380 120880 123620 120900
rect 123880 120880 124120 120900
rect 124380 120880 124620 120900
rect 124880 120880 125120 120900
rect 125380 120880 125620 120900
rect 125880 120880 126120 120900
rect 126380 120880 126620 120900
rect 126880 120880 127120 120900
rect 127380 120880 127620 120900
rect 127880 120880 128120 120900
rect 128380 120880 128620 120900
rect 128880 120880 129120 120900
rect 129380 120880 129620 120900
rect 129880 120880 130120 120900
rect 130380 120880 130620 120900
rect 130880 120880 131120 120900
rect 131380 120880 131620 120900
rect 131880 120880 132120 120900
rect 132380 120880 132620 120900
rect 132880 120880 133120 120900
rect 133380 120880 133620 120900
rect 133880 120880 134120 120900
rect 134380 120880 134620 120900
rect 134880 120880 135120 120900
rect 135380 120880 135620 120900
rect 135880 120880 136120 120900
rect 136380 120880 136620 120900
rect 136880 120880 137120 120900
rect 137380 120880 137620 120900
rect 137880 120880 138120 120900
rect 138380 120880 138620 120900
rect 138880 120880 139120 120900
rect 139380 120880 139620 120900
rect 139880 120880 140120 120900
rect 140380 120880 140620 120900
rect 140880 120880 141120 120900
rect 141380 120880 141620 120900
rect 141880 120880 142000 120900
rect 118000 120620 118100 120880
rect 118400 120620 118600 120880
rect 118900 120620 119100 120880
rect 119400 120620 119600 120880
rect 119900 120620 120100 120880
rect 120400 120620 120600 120880
rect 120900 120620 121100 120880
rect 121400 120620 121600 120880
rect 121900 120620 122100 120880
rect 122400 120620 122600 120880
rect 122900 120620 123100 120880
rect 123400 120620 123600 120880
rect 123900 120620 124100 120880
rect 124400 120620 124600 120880
rect 124900 120620 125100 120880
rect 125400 120620 125600 120880
rect 125900 120620 126100 120880
rect 126400 120620 126600 120880
rect 126900 120620 127100 120880
rect 127400 120620 127600 120880
rect 127900 120620 128100 120880
rect 128400 120620 128600 120880
rect 128900 120620 129100 120880
rect 129400 120620 129600 120880
rect 129900 120620 130100 120880
rect 130400 120620 130600 120880
rect 130900 120620 131100 120880
rect 131400 120620 131600 120880
rect 131900 120620 132100 120880
rect 132400 120620 132600 120880
rect 132900 120620 133100 120880
rect 133400 120620 133600 120880
rect 133900 120620 134100 120880
rect 134400 120620 134600 120880
rect 134900 120620 135100 120880
rect 135400 120620 135600 120880
rect 135900 120620 136100 120880
rect 136400 120620 136600 120880
rect 136900 120620 137100 120880
rect 137400 120620 137600 120880
rect 137900 120620 138100 120880
rect 138400 120620 138600 120880
rect 138900 120620 139100 120880
rect 139400 120620 139600 120880
rect 139900 120620 140100 120880
rect 140400 120620 140600 120880
rect 140900 120620 141100 120880
rect 141400 120620 141600 120880
rect 141900 120620 142000 120880
rect 118000 120600 118120 120620
rect 118380 120600 118620 120620
rect 118880 120600 119120 120620
rect 119380 120600 119620 120620
rect 119880 120600 120120 120620
rect 120380 120600 120620 120620
rect 120880 120600 121120 120620
rect 121380 120600 121620 120620
rect 121880 120600 122120 120620
rect 122380 120600 122620 120620
rect 122880 120600 123120 120620
rect 123380 120600 123620 120620
rect 123880 120600 124120 120620
rect 124380 120600 124620 120620
rect 124880 120600 125120 120620
rect 125380 120600 125620 120620
rect 125880 120600 126120 120620
rect 126380 120600 126620 120620
rect 126880 120600 127120 120620
rect 127380 120600 127620 120620
rect 127880 120600 128120 120620
rect 128380 120600 128620 120620
rect 128880 120600 129120 120620
rect 129380 120600 129620 120620
rect 129880 120600 130120 120620
rect 130380 120600 130620 120620
rect 130880 120600 131120 120620
rect 131380 120600 131620 120620
rect 131880 120600 132120 120620
rect 132380 120600 132620 120620
rect 132880 120600 133120 120620
rect 133380 120600 133620 120620
rect 133880 120600 134120 120620
rect 134380 120600 134620 120620
rect 134880 120600 135120 120620
rect 135380 120600 135620 120620
rect 135880 120600 136120 120620
rect 136380 120600 136620 120620
rect 136880 120600 137120 120620
rect 137380 120600 137620 120620
rect 137880 120600 138120 120620
rect 138380 120600 138620 120620
rect 138880 120600 139120 120620
rect 139380 120600 139620 120620
rect 139880 120600 140120 120620
rect 140380 120600 140620 120620
rect 140880 120600 141120 120620
rect 141380 120600 141620 120620
rect 141880 120600 142000 120620
rect 118000 120400 142000 120600
rect 118000 120380 118120 120400
rect 118380 120380 118620 120400
rect 118880 120380 119120 120400
rect 119380 120380 119620 120400
rect 119880 120380 120120 120400
rect 120380 120380 120620 120400
rect 120880 120380 121120 120400
rect 121380 120380 121620 120400
rect 121880 120380 122120 120400
rect 122380 120380 122620 120400
rect 122880 120380 123120 120400
rect 123380 120380 123620 120400
rect 123880 120380 124120 120400
rect 124380 120380 124620 120400
rect 124880 120380 125120 120400
rect 125380 120380 125620 120400
rect 125880 120380 126120 120400
rect 126380 120380 126620 120400
rect 126880 120380 127120 120400
rect 127380 120380 127620 120400
rect 127880 120380 128120 120400
rect 128380 120380 128620 120400
rect 128880 120380 129120 120400
rect 129380 120380 129620 120400
rect 129880 120380 130120 120400
rect 130380 120380 130620 120400
rect 130880 120380 131120 120400
rect 131380 120380 131620 120400
rect 131880 120380 132120 120400
rect 132380 120380 132620 120400
rect 132880 120380 133120 120400
rect 133380 120380 133620 120400
rect 133880 120380 134120 120400
rect 134380 120380 134620 120400
rect 134880 120380 135120 120400
rect 135380 120380 135620 120400
rect 135880 120380 136120 120400
rect 136380 120380 136620 120400
rect 136880 120380 137120 120400
rect 137380 120380 137620 120400
rect 137880 120380 138120 120400
rect 138380 120380 138620 120400
rect 138880 120380 139120 120400
rect 139380 120380 139620 120400
rect 139880 120380 140120 120400
rect 140380 120380 140620 120400
rect 140880 120380 141120 120400
rect 141380 120380 141620 120400
rect 141880 120380 142000 120400
rect 118000 120120 118100 120380
rect 118400 120120 118600 120380
rect 118900 120120 119100 120380
rect 119400 120120 119600 120380
rect 119900 120120 120100 120380
rect 120400 120120 120600 120380
rect 120900 120120 121100 120380
rect 121400 120120 121600 120380
rect 121900 120120 122100 120380
rect 122400 120120 122600 120380
rect 122900 120120 123100 120380
rect 123400 120120 123600 120380
rect 123900 120120 124100 120380
rect 124400 120120 124600 120380
rect 124900 120120 125100 120380
rect 125400 120120 125600 120380
rect 125900 120120 126100 120380
rect 126400 120120 126600 120380
rect 126900 120120 127100 120380
rect 127400 120120 127600 120380
rect 127900 120120 128100 120380
rect 128400 120120 128600 120380
rect 128900 120120 129100 120380
rect 129400 120120 129600 120380
rect 129900 120120 130100 120380
rect 130400 120120 130600 120380
rect 130900 120120 131100 120380
rect 131400 120120 131600 120380
rect 131900 120120 132100 120380
rect 132400 120120 132600 120380
rect 132900 120120 133100 120380
rect 133400 120120 133600 120380
rect 133900 120120 134100 120380
rect 134400 120120 134600 120380
rect 134900 120120 135100 120380
rect 135400 120120 135600 120380
rect 135900 120120 136100 120380
rect 136400 120120 136600 120380
rect 136900 120120 137100 120380
rect 137400 120120 137600 120380
rect 137900 120120 138100 120380
rect 138400 120120 138600 120380
rect 138900 120120 139100 120380
rect 139400 120120 139600 120380
rect 139900 120120 140100 120380
rect 140400 120120 140600 120380
rect 140900 120120 141100 120380
rect 141400 120120 141600 120380
rect 141900 120120 142000 120380
rect 118000 120100 118120 120120
rect 118380 120100 118620 120120
rect 118880 120100 119120 120120
rect 119380 120100 119620 120120
rect 119880 120100 120120 120120
rect 120380 120100 120620 120120
rect 120880 120100 121120 120120
rect 121380 120100 121620 120120
rect 121880 120100 122120 120120
rect 122380 120100 122620 120120
rect 122880 120100 123120 120120
rect 123380 120100 123620 120120
rect 123880 120100 124120 120120
rect 124380 120100 124620 120120
rect 124880 120100 125120 120120
rect 125380 120100 125620 120120
rect 125880 120100 126120 120120
rect 126380 120100 126620 120120
rect 126880 120100 127120 120120
rect 127380 120100 127620 120120
rect 127880 120100 128120 120120
rect 128380 120100 128620 120120
rect 128880 120100 129120 120120
rect 129380 120100 129620 120120
rect 129880 120100 130120 120120
rect 130380 120100 130620 120120
rect 130880 120100 131120 120120
rect 131380 120100 131620 120120
rect 131880 120100 132120 120120
rect 132380 120100 132620 120120
rect 132880 120100 133120 120120
rect 133380 120100 133620 120120
rect 133880 120100 134120 120120
rect 134380 120100 134620 120120
rect 134880 120100 135120 120120
rect 135380 120100 135620 120120
rect 135880 120100 136120 120120
rect 136380 120100 136620 120120
rect 136880 120100 137120 120120
rect 137380 120100 137620 120120
rect 137880 120100 138120 120120
rect 138380 120100 138620 120120
rect 138880 120100 139120 120120
rect 139380 120100 139620 120120
rect 139880 120100 140120 120120
rect 140380 120100 140620 120120
rect 140880 120100 141120 120120
rect 141380 120100 141620 120120
rect 141880 120100 142000 120120
rect 118000 119900 142000 120100
rect 118000 119880 118120 119900
rect 118380 119880 118620 119900
rect 118880 119880 119120 119900
rect 119380 119880 119620 119900
rect 119880 119880 120120 119900
rect 120380 119880 120620 119900
rect 120880 119880 121120 119900
rect 121380 119880 121620 119900
rect 121880 119880 122120 119900
rect 122380 119880 122620 119900
rect 122880 119880 123120 119900
rect 123380 119880 123620 119900
rect 123880 119880 124120 119900
rect 124380 119880 124620 119900
rect 124880 119880 125120 119900
rect 125380 119880 125620 119900
rect 125880 119880 126120 119900
rect 126380 119880 126620 119900
rect 126880 119880 127120 119900
rect 127380 119880 127620 119900
rect 127880 119880 128120 119900
rect 128380 119880 128620 119900
rect 128880 119880 129120 119900
rect 129380 119880 129620 119900
rect 129880 119880 130120 119900
rect 130380 119880 130620 119900
rect 130880 119880 131120 119900
rect 131380 119880 131620 119900
rect 131880 119880 132120 119900
rect 132380 119880 132620 119900
rect 132880 119880 133120 119900
rect 133380 119880 133620 119900
rect 133880 119880 134120 119900
rect 134380 119880 134620 119900
rect 134880 119880 135120 119900
rect 135380 119880 135620 119900
rect 135880 119880 136120 119900
rect 136380 119880 136620 119900
rect 136880 119880 137120 119900
rect 137380 119880 137620 119900
rect 137880 119880 138120 119900
rect 138380 119880 138620 119900
rect 138880 119880 139120 119900
rect 139380 119880 139620 119900
rect 139880 119880 140120 119900
rect 140380 119880 140620 119900
rect 140880 119880 141120 119900
rect 141380 119880 141620 119900
rect 141880 119880 142000 119900
rect 118000 119620 118100 119880
rect 118400 119620 118600 119880
rect 118900 119620 119100 119880
rect 119400 119620 119600 119880
rect 119900 119620 120100 119880
rect 120400 119620 120600 119880
rect 120900 119620 121100 119880
rect 121400 119620 121600 119880
rect 121900 119620 122100 119880
rect 122400 119620 122600 119880
rect 122900 119620 123100 119880
rect 123400 119620 123600 119880
rect 123900 119620 124100 119880
rect 124400 119620 124600 119880
rect 124900 119620 125100 119880
rect 125400 119620 125600 119880
rect 125900 119620 126100 119880
rect 126400 119620 126600 119880
rect 126900 119620 127100 119880
rect 127400 119620 127600 119880
rect 127900 119620 128100 119880
rect 128400 119620 128600 119880
rect 128900 119620 129100 119880
rect 129400 119620 129600 119880
rect 129900 119620 130100 119880
rect 130400 119620 130600 119880
rect 130900 119620 131100 119880
rect 131400 119620 131600 119880
rect 131900 119620 132100 119880
rect 132400 119620 132600 119880
rect 132900 119620 133100 119880
rect 133400 119620 133600 119880
rect 133900 119620 134100 119880
rect 134400 119620 134600 119880
rect 134900 119620 135100 119880
rect 135400 119620 135600 119880
rect 135900 119620 136100 119880
rect 136400 119620 136600 119880
rect 136900 119620 137100 119880
rect 137400 119620 137600 119880
rect 137900 119620 138100 119880
rect 138400 119620 138600 119880
rect 138900 119620 139100 119880
rect 139400 119620 139600 119880
rect 139900 119620 140100 119880
rect 140400 119620 140600 119880
rect 140900 119620 141100 119880
rect 141400 119620 141600 119880
rect 141900 119620 142000 119880
rect 118000 119600 118120 119620
rect 118380 119600 118620 119620
rect 118880 119600 119120 119620
rect 119380 119600 119620 119620
rect 119880 119600 120120 119620
rect 120380 119600 120620 119620
rect 120880 119600 121120 119620
rect 121380 119600 121620 119620
rect 121880 119600 122120 119620
rect 122380 119600 122620 119620
rect 122880 119600 123120 119620
rect 123380 119600 123620 119620
rect 123880 119600 124120 119620
rect 124380 119600 124620 119620
rect 124880 119600 125120 119620
rect 125380 119600 125620 119620
rect 125880 119600 126120 119620
rect 126380 119600 126620 119620
rect 126880 119600 127120 119620
rect 127380 119600 127620 119620
rect 127880 119600 128120 119620
rect 128380 119600 128620 119620
rect 128880 119600 129120 119620
rect 129380 119600 129620 119620
rect 129880 119600 130120 119620
rect 130380 119600 130620 119620
rect 130880 119600 131120 119620
rect 131380 119600 131620 119620
rect 131880 119600 132120 119620
rect 132380 119600 132620 119620
rect 132880 119600 133120 119620
rect 133380 119600 133620 119620
rect 133880 119600 134120 119620
rect 134380 119600 134620 119620
rect 134880 119600 135120 119620
rect 135380 119600 135620 119620
rect 135880 119600 136120 119620
rect 136380 119600 136620 119620
rect 136880 119600 137120 119620
rect 137380 119600 137620 119620
rect 137880 119600 138120 119620
rect 138380 119600 138620 119620
rect 138880 119600 139120 119620
rect 139380 119600 139620 119620
rect 139880 119600 140120 119620
rect 140380 119600 140620 119620
rect 140880 119600 141120 119620
rect 141380 119600 141620 119620
rect 141880 119600 142000 119620
rect 118000 119400 142000 119600
rect 118000 119380 118120 119400
rect 118380 119380 118620 119400
rect 118880 119380 119120 119400
rect 119380 119380 119620 119400
rect 119880 119380 120120 119400
rect 120380 119380 120620 119400
rect 120880 119380 121120 119400
rect 121380 119380 121620 119400
rect 121880 119380 122120 119400
rect 122380 119380 122620 119400
rect 122880 119380 123120 119400
rect 123380 119380 123620 119400
rect 123880 119380 124120 119400
rect 124380 119380 124620 119400
rect 124880 119380 125120 119400
rect 125380 119380 125620 119400
rect 125880 119380 126120 119400
rect 126380 119380 126620 119400
rect 126880 119380 127120 119400
rect 127380 119380 127620 119400
rect 127880 119380 128120 119400
rect 128380 119380 128620 119400
rect 128880 119380 129120 119400
rect 129380 119380 129620 119400
rect 129880 119380 130120 119400
rect 130380 119380 130620 119400
rect 130880 119380 131120 119400
rect 131380 119380 131620 119400
rect 131880 119380 132120 119400
rect 132380 119380 132620 119400
rect 132880 119380 133120 119400
rect 133380 119380 133620 119400
rect 133880 119380 134120 119400
rect 134380 119380 134620 119400
rect 134880 119380 135120 119400
rect 135380 119380 135620 119400
rect 135880 119380 136120 119400
rect 136380 119380 136620 119400
rect 136880 119380 137120 119400
rect 137380 119380 137620 119400
rect 137880 119380 138120 119400
rect 138380 119380 138620 119400
rect 138880 119380 139120 119400
rect 139380 119380 139620 119400
rect 139880 119380 140120 119400
rect 140380 119380 140620 119400
rect 140880 119380 141120 119400
rect 141380 119380 141620 119400
rect 141880 119380 142000 119400
rect 118000 119120 118100 119380
rect 118400 119120 118600 119380
rect 118900 119120 119100 119380
rect 119400 119120 119600 119380
rect 119900 119120 120100 119380
rect 120400 119120 120600 119380
rect 120900 119120 121100 119380
rect 121400 119120 121600 119380
rect 121900 119120 122100 119380
rect 122400 119120 122600 119380
rect 122900 119120 123100 119380
rect 123400 119120 123600 119380
rect 123900 119120 124100 119380
rect 124400 119120 124600 119380
rect 124900 119120 125100 119380
rect 125400 119120 125600 119380
rect 125900 119120 126100 119380
rect 126400 119120 126600 119380
rect 126900 119120 127100 119380
rect 127400 119120 127600 119380
rect 127900 119120 128100 119380
rect 128400 119120 128600 119380
rect 128900 119120 129100 119380
rect 129400 119120 129600 119380
rect 129900 119120 130100 119380
rect 130400 119120 130600 119380
rect 130900 119120 131100 119380
rect 131400 119120 131600 119380
rect 131900 119120 132100 119380
rect 132400 119120 132600 119380
rect 132900 119120 133100 119380
rect 133400 119120 133600 119380
rect 133900 119120 134100 119380
rect 134400 119120 134600 119380
rect 134900 119120 135100 119380
rect 135400 119120 135600 119380
rect 135900 119120 136100 119380
rect 136400 119120 136600 119380
rect 136900 119120 137100 119380
rect 137400 119120 137600 119380
rect 137900 119120 138100 119380
rect 138400 119120 138600 119380
rect 138900 119120 139100 119380
rect 139400 119120 139600 119380
rect 139900 119120 140100 119380
rect 140400 119120 140600 119380
rect 140900 119120 141100 119380
rect 141400 119120 141600 119380
rect 141900 119120 142000 119380
rect 118000 119100 118120 119120
rect 118380 119100 118620 119120
rect 118880 119100 119120 119120
rect 119380 119100 119620 119120
rect 119880 119100 120120 119120
rect 120380 119100 120620 119120
rect 120880 119100 121120 119120
rect 121380 119100 121620 119120
rect 121880 119100 122120 119120
rect 122380 119100 122620 119120
rect 122880 119100 123120 119120
rect 123380 119100 123620 119120
rect 123880 119100 124120 119120
rect 124380 119100 124620 119120
rect 124880 119100 125120 119120
rect 125380 119100 125620 119120
rect 125880 119100 126120 119120
rect 126380 119100 126620 119120
rect 126880 119100 127120 119120
rect 127380 119100 127620 119120
rect 127880 119100 128120 119120
rect 128380 119100 128620 119120
rect 128880 119100 129120 119120
rect 129380 119100 129620 119120
rect 129880 119100 130120 119120
rect 130380 119100 130620 119120
rect 130880 119100 131120 119120
rect 131380 119100 131620 119120
rect 131880 119100 132120 119120
rect 132380 119100 132620 119120
rect 132880 119100 133120 119120
rect 133380 119100 133620 119120
rect 133880 119100 134120 119120
rect 134380 119100 134620 119120
rect 134880 119100 135120 119120
rect 135380 119100 135620 119120
rect 135880 119100 136120 119120
rect 136380 119100 136620 119120
rect 136880 119100 137120 119120
rect 137380 119100 137620 119120
rect 137880 119100 138120 119120
rect 138380 119100 138620 119120
rect 138880 119100 139120 119120
rect 139380 119100 139620 119120
rect 139880 119100 140120 119120
rect 140380 119100 140620 119120
rect 140880 119100 141120 119120
rect 141380 119100 141620 119120
rect 141880 119100 142000 119120
rect 118000 118900 142000 119100
rect 118000 118880 118120 118900
rect 118380 118880 118620 118900
rect 118880 118880 119120 118900
rect 119380 118880 119620 118900
rect 119880 118880 120120 118900
rect 120380 118880 120620 118900
rect 120880 118880 121120 118900
rect 121380 118880 121620 118900
rect 121880 118880 122120 118900
rect 122380 118880 122620 118900
rect 122880 118880 123120 118900
rect 123380 118880 123620 118900
rect 123880 118880 124120 118900
rect 124380 118880 124620 118900
rect 124880 118880 125120 118900
rect 125380 118880 125620 118900
rect 125880 118880 126120 118900
rect 126380 118880 126620 118900
rect 126880 118880 127120 118900
rect 127380 118880 127620 118900
rect 127880 118880 128120 118900
rect 128380 118880 128620 118900
rect 128880 118880 129120 118900
rect 129380 118880 129620 118900
rect 129880 118880 130120 118900
rect 130380 118880 130620 118900
rect 130880 118880 131120 118900
rect 131380 118880 131620 118900
rect 131880 118880 132120 118900
rect 132380 118880 132620 118900
rect 132880 118880 133120 118900
rect 133380 118880 133620 118900
rect 133880 118880 134120 118900
rect 134380 118880 134620 118900
rect 134880 118880 135120 118900
rect 135380 118880 135620 118900
rect 135880 118880 136120 118900
rect 136380 118880 136620 118900
rect 136880 118880 137120 118900
rect 137380 118880 137620 118900
rect 137880 118880 138120 118900
rect 138380 118880 138620 118900
rect 138880 118880 139120 118900
rect 139380 118880 139620 118900
rect 139880 118880 140120 118900
rect 140380 118880 140620 118900
rect 140880 118880 141120 118900
rect 141380 118880 141620 118900
rect 141880 118880 142000 118900
rect 118000 118620 118100 118880
rect 118400 118620 118600 118880
rect 118900 118620 119100 118880
rect 119400 118620 119600 118880
rect 119900 118620 120100 118880
rect 120400 118620 120600 118880
rect 120900 118620 121100 118880
rect 121400 118620 121600 118880
rect 121900 118620 122100 118880
rect 122400 118620 122600 118880
rect 122900 118620 123100 118880
rect 123400 118620 123600 118880
rect 123900 118620 124100 118880
rect 124400 118620 124600 118880
rect 124900 118620 125100 118880
rect 125400 118620 125600 118880
rect 125900 118620 126100 118880
rect 126400 118620 126600 118880
rect 126900 118620 127100 118880
rect 127400 118620 127600 118880
rect 127900 118620 128100 118880
rect 128400 118620 128600 118880
rect 128900 118620 129100 118880
rect 129400 118620 129600 118880
rect 129900 118620 130100 118880
rect 130400 118620 130600 118880
rect 130900 118620 131100 118880
rect 131400 118620 131600 118880
rect 131900 118620 132100 118880
rect 132400 118620 132600 118880
rect 132900 118620 133100 118880
rect 133400 118620 133600 118880
rect 133900 118620 134100 118880
rect 134400 118620 134600 118880
rect 134900 118620 135100 118880
rect 135400 118620 135600 118880
rect 135900 118620 136100 118880
rect 136400 118620 136600 118880
rect 136900 118620 137100 118880
rect 137400 118620 137600 118880
rect 137900 118620 138100 118880
rect 138400 118620 138600 118880
rect 138900 118620 139100 118880
rect 139400 118620 139600 118880
rect 139900 118620 140100 118880
rect 140400 118620 140600 118880
rect 140900 118620 141100 118880
rect 141400 118620 141600 118880
rect 141900 118620 142000 118880
rect 118000 118600 118120 118620
rect 118380 118600 118620 118620
rect 118880 118600 119120 118620
rect 119380 118600 119620 118620
rect 119880 118600 120120 118620
rect 120380 118600 120620 118620
rect 120880 118600 121120 118620
rect 121380 118600 121620 118620
rect 121880 118600 122120 118620
rect 122380 118600 122620 118620
rect 122880 118600 123120 118620
rect 123380 118600 123620 118620
rect 123880 118600 124120 118620
rect 124380 118600 124620 118620
rect 124880 118600 125120 118620
rect 125380 118600 125620 118620
rect 125880 118600 126120 118620
rect 126380 118600 126620 118620
rect 126880 118600 127120 118620
rect 127380 118600 127620 118620
rect 127880 118600 128120 118620
rect 128380 118600 128620 118620
rect 128880 118600 129120 118620
rect 129380 118600 129620 118620
rect 129880 118600 130120 118620
rect 130380 118600 130620 118620
rect 130880 118600 131120 118620
rect 131380 118600 131620 118620
rect 131880 118600 132120 118620
rect 132380 118600 132620 118620
rect 132880 118600 133120 118620
rect 133380 118600 133620 118620
rect 133880 118600 134120 118620
rect 134380 118600 134620 118620
rect 134880 118600 135120 118620
rect 135380 118600 135620 118620
rect 135880 118600 136120 118620
rect 136380 118600 136620 118620
rect 136880 118600 137120 118620
rect 137380 118600 137620 118620
rect 137880 118600 138120 118620
rect 138380 118600 138620 118620
rect 138880 118600 139120 118620
rect 139380 118600 139620 118620
rect 139880 118600 140120 118620
rect 140380 118600 140620 118620
rect 140880 118600 141120 118620
rect 141380 118600 141620 118620
rect 141880 118600 142000 118620
rect 118000 118400 142000 118600
rect 118000 118380 118120 118400
rect 118380 118380 118620 118400
rect 118880 118380 119120 118400
rect 119380 118380 119620 118400
rect 119880 118380 120120 118400
rect 120380 118380 120620 118400
rect 120880 118380 121120 118400
rect 121380 118380 121620 118400
rect 121880 118380 122120 118400
rect 122380 118380 122620 118400
rect 122880 118380 123120 118400
rect 123380 118380 123620 118400
rect 123880 118380 124120 118400
rect 124380 118380 124620 118400
rect 124880 118380 125120 118400
rect 125380 118380 125620 118400
rect 125880 118380 126120 118400
rect 126380 118380 126620 118400
rect 126880 118380 127120 118400
rect 127380 118380 127620 118400
rect 127880 118380 128120 118400
rect 128380 118380 128620 118400
rect 128880 118380 129120 118400
rect 129380 118380 129620 118400
rect 129880 118380 130120 118400
rect 130380 118380 130620 118400
rect 130880 118380 131120 118400
rect 131380 118380 131620 118400
rect 131880 118380 132120 118400
rect 132380 118380 132620 118400
rect 132880 118380 133120 118400
rect 133380 118380 133620 118400
rect 133880 118380 134120 118400
rect 134380 118380 134620 118400
rect 134880 118380 135120 118400
rect 135380 118380 135620 118400
rect 135880 118380 136120 118400
rect 136380 118380 136620 118400
rect 136880 118380 137120 118400
rect 137380 118380 137620 118400
rect 137880 118380 138120 118400
rect 138380 118380 138620 118400
rect 138880 118380 139120 118400
rect 139380 118380 139620 118400
rect 139880 118380 140120 118400
rect 140380 118380 140620 118400
rect 140880 118380 141120 118400
rect 141380 118380 141620 118400
rect 141880 118380 142000 118400
rect 118000 118120 118100 118380
rect 118400 118120 118600 118380
rect 118900 118120 119100 118380
rect 119400 118120 119600 118380
rect 119900 118120 120100 118380
rect 120400 118120 120600 118380
rect 120900 118120 121100 118380
rect 121400 118120 121600 118380
rect 121900 118120 122100 118380
rect 122400 118120 122600 118380
rect 122900 118120 123100 118380
rect 123400 118120 123600 118380
rect 123900 118120 124100 118380
rect 124400 118120 124600 118380
rect 124900 118120 125100 118380
rect 125400 118120 125600 118380
rect 125900 118120 126100 118380
rect 126400 118120 126600 118380
rect 126900 118120 127100 118380
rect 127400 118120 127600 118380
rect 127900 118120 128100 118380
rect 128400 118120 128600 118380
rect 128900 118120 129100 118380
rect 129400 118120 129600 118380
rect 129900 118120 130100 118380
rect 130400 118120 130600 118380
rect 130900 118120 131100 118380
rect 131400 118120 131600 118380
rect 131900 118120 132100 118380
rect 132400 118120 132600 118380
rect 132900 118120 133100 118380
rect 133400 118120 133600 118380
rect 133900 118120 134100 118380
rect 134400 118120 134600 118380
rect 134900 118120 135100 118380
rect 135400 118120 135600 118380
rect 135900 118120 136100 118380
rect 136400 118120 136600 118380
rect 136900 118120 137100 118380
rect 137400 118120 137600 118380
rect 137900 118120 138100 118380
rect 138400 118120 138600 118380
rect 138900 118120 139100 118380
rect 139400 118120 139600 118380
rect 139900 118120 140100 118380
rect 140400 118120 140600 118380
rect 140900 118120 141100 118380
rect 141400 118120 141600 118380
rect 141900 118120 142000 118380
rect 118000 118100 118120 118120
rect 118380 118100 118620 118120
rect 118880 118100 119120 118120
rect 119380 118100 119620 118120
rect 119880 118100 120120 118120
rect 120380 118100 120620 118120
rect 120880 118100 121120 118120
rect 121380 118100 121620 118120
rect 121880 118100 122120 118120
rect 122380 118100 122620 118120
rect 122880 118100 123120 118120
rect 123380 118100 123620 118120
rect 123880 118100 124120 118120
rect 124380 118100 124620 118120
rect 124880 118100 125120 118120
rect 125380 118100 125620 118120
rect 125880 118100 126120 118120
rect 126380 118100 126620 118120
rect 126880 118100 127120 118120
rect 127380 118100 127620 118120
rect 127880 118100 128120 118120
rect 128380 118100 128620 118120
rect 128880 118100 129120 118120
rect 129380 118100 129620 118120
rect 129880 118100 130120 118120
rect 130380 118100 130620 118120
rect 130880 118100 131120 118120
rect 131380 118100 131620 118120
rect 131880 118100 132120 118120
rect 132380 118100 132620 118120
rect 132880 118100 133120 118120
rect 133380 118100 133620 118120
rect 133880 118100 134120 118120
rect 134380 118100 134620 118120
rect 134880 118100 135120 118120
rect 135380 118100 135620 118120
rect 135880 118100 136120 118120
rect 136380 118100 136620 118120
rect 136880 118100 137120 118120
rect 137380 118100 137620 118120
rect 137880 118100 138120 118120
rect 138380 118100 138620 118120
rect 138880 118100 139120 118120
rect 139380 118100 139620 118120
rect 139880 118100 140120 118120
rect 140380 118100 140620 118120
rect 140880 118100 141120 118120
rect 141380 118100 141620 118120
rect 141880 118100 142000 118120
rect 118000 117900 142000 118100
rect 118000 117880 118120 117900
rect 118380 117880 118620 117900
rect 118880 117880 119120 117900
rect 119380 117880 119620 117900
rect 119880 117880 120120 117900
rect 120380 117880 120620 117900
rect 120880 117880 121120 117900
rect 121380 117880 121620 117900
rect 121880 117880 122120 117900
rect 122380 117880 122620 117900
rect 122880 117880 123120 117900
rect 123380 117880 123620 117900
rect 123880 117880 124120 117900
rect 124380 117880 124620 117900
rect 124880 117880 125120 117900
rect 125380 117880 125620 117900
rect 125880 117880 126120 117900
rect 126380 117880 126620 117900
rect 126880 117880 127120 117900
rect 127380 117880 127620 117900
rect 127880 117880 128120 117900
rect 128380 117880 128620 117900
rect 128880 117880 129120 117900
rect 129380 117880 129620 117900
rect 129880 117880 130120 117900
rect 130380 117880 130620 117900
rect 130880 117880 131120 117900
rect 131380 117880 131620 117900
rect 131880 117880 132120 117900
rect 132380 117880 132620 117900
rect 132880 117880 133120 117900
rect 133380 117880 133620 117900
rect 133880 117880 134120 117900
rect 134380 117880 134620 117900
rect 134880 117880 135120 117900
rect 135380 117880 135620 117900
rect 135880 117880 136120 117900
rect 136380 117880 136620 117900
rect 136880 117880 137120 117900
rect 137380 117880 137620 117900
rect 137880 117880 138120 117900
rect 138380 117880 138620 117900
rect 138880 117880 139120 117900
rect 139380 117880 139620 117900
rect 139880 117880 140120 117900
rect 140380 117880 140620 117900
rect 140880 117880 141120 117900
rect 141380 117880 141620 117900
rect 141880 117880 142000 117900
rect 118000 117620 118100 117880
rect 118400 117620 118600 117880
rect 118900 117620 119100 117880
rect 119400 117620 119600 117880
rect 119900 117620 120100 117880
rect 120400 117620 120600 117880
rect 120900 117620 121100 117880
rect 121400 117620 121600 117880
rect 121900 117620 122100 117880
rect 122400 117620 122600 117880
rect 122900 117620 123100 117880
rect 123400 117620 123600 117880
rect 123900 117620 124100 117880
rect 124400 117620 124600 117880
rect 124900 117620 125100 117880
rect 125400 117620 125600 117880
rect 125900 117620 126100 117880
rect 126400 117620 126600 117880
rect 126900 117620 127100 117880
rect 127400 117620 127600 117880
rect 127900 117620 128100 117880
rect 128400 117620 128600 117880
rect 128900 117620 129100 117880
rect 129400 117620 129600 117880
rect 129900 117620 130100 117880
rect 130400 117620 130600 117880
rect 130900 117620 131100 117880
rect 131400 117620 131600 117880
rect 131900 117620 132100 117880
rect 132400 117620 132600 117880
rect 132900 117620 133100 117880
rect 133400 117620 133600 117880
rect 133900 117620 134100 117880
rect 134400 117620 134600 117880
rect 134900 117620 135100 117880
rect 135400 117620 135600 117880
rect 135900 117620 136100 117880
rect 136400 117620 136600 117880
rect 136900 117620 137100 117880
rect 137400 117620 137600 117880
rect 137900 117620 138100 117880
rect 138400 117620 138600 117880
rect 138900 117620 139100 117880
rect 139400 117620 139600 117880
rect 139900 117620 140100 117880
rect 140400 117620 140600 117880
rect 140900 117620 141100 117880
rect 141400 117620 141600 117880
rect 141900 117620 142000 117880
rect 118000 117600 118120 117620
rect 118380 117600 118620 117620
rect 118880 117600 119120 117620
rect 119380 117600 119620 117620
rect 119880 117600 120120 117620
rect 120380 117600 120620 117620
rect 120880 117600 121120 117620
rect 121380 117600 121620 117620
rect 121880 117600 122120 117620
rect 122380 117600 122620 117620
rect 122880 117600 123120 117620
rect 123380 117600 123620 117620
rect 123880 117600 124120 117620
rect 124380 117600 124620 117620
rect 124880 117600 125120 117620
rect 125380 117600 125620 117620
rect 125880 117600 126120 117620
rect 126380 117600 126620 117620
rect 126880 117600 127120 117620
rect 127380 117600 127620 117620
rect 127880 117600 128120 117620
rect 128380 117600 128620 117620
rect 128880 117600 129120 117620
rect 129380 117600 129620 117620
rect 129880 117600 130120 117620
rect 130380 117600 130620 117620
rect 130880 117600 131120 117620
rect 131380 117600 131620 117620
rect 131880 117600 132120 117620
rect 132380 117600 132620 117620
rect 132880 117600 133120 117620
rect 133380 117600 133620 117620
rect 133880 117600 134120 117620
rect 134380 117600 134620 117620
rect 134880 117600 135120 117620
rect 135380 117600 135620 117620
rect 135880 117600 136120 117620
rect 136380 117600 136620 117620
rect 136880 117600 137120 117620
rect 137380 117600 137620 117620
rect 137880 117600 138120 117620
rect 138380 117600 138620 117620
rect 138880 117600 139120 117620
rect 139380 117600 139620 117620
rect 139880 117600 140120 117620
rect 140380 117600 140620 117620
rect 140880 117600 141120 117620
rect 141380 117600 141620 117620
rect 141880 117600 142000 117620
rect 118000 117400 142000 117600
rect 118000 117380 118120 117400
rect 118380 117380 118620 117400
rect 118880 117380 119120 117400
rect 119380 117380 119620 117400
rect 119880 117380 120120 117400
rect 120380 117380 120620 117400
rect 120880 117380 121120 117400
rect 121380 117380 121620 117400
rect 121880 117380 122120 117400
rect 122380 117380 122620 117400
rect 122880 117380 123120 117400
rect 123380 117380 123620 117400
rect 123880 117380 124120 117400
rect 124380 117380 124620 117400
rect 124880 117380 125120 117400
rect 125380 117380 125620 117400
rect 125880 117380 126120 117400
rect 126380 117380 126620 117400
rect 126880 117380 127120 117400
rect 127380 117380 127620 117400
rect 127880 117380 128120 117400
rect 128380 117380 128620 117400
rect 128880 117380 129120 117400
rect 129380 117380 129620 117400
rect 129880 117380 130120 117400
rect 130380 117380 130620 117400
rect 130880 117380 131120 117400
rect 131380 117380 131620 117400
rect 131880 117380 132120 117400
rect 132380 117380 132620 117400
rect 132880 117380 133120 117400
rect 133380 117380 133620 117400
rect 133880 117380 134120 117400
rect 134380 117380 134620 117400
rect 134880 117380 135120 117400
rect 135380 117380 135620 117400
rect 135880 117380 136120 117400
rect 136380 117380 136620 117400
rect 136880 117380 137120 117400
rect 137380 117380 137620 117400
rect 137880 117380 138120 117400
rect 138380 117380 138620 117400
rect 138880 117380 139120 117400
rect 139380 117380 139620 117400
rect 139880 117380 140120 117400
rect 140380 117380 140620 117400
rect 140880 117380 141120 117400
rect 141380 117380 141620 117400
rect 141880 117380 142000 117400
rect 118000 117120 118100 117380
rect 118400 117120 118600 117380
rect 118900 117120 119100 117380
rect 119400 117120 119600 117380
rect 119900 117120 120100 117380
rect 120400 117120 120600 117380
rect 120900 117120 121100 117380
rect 121400 117120 121600 117380
rect 121900 117120 122100 117380
rect 122400 117120 122600 117380
rect 122900 117120 123100 117380
rect 123400 117120 123600 117380
rect 123900 117120 124100 117380
rect 124400 117120 124600 117380
rect 124900 117120 125100 117380
rect 125400 117120 125600 117380
rect 125900 117120 126100 117380
rect 126400 117120 126600 117380
rect 126900 117120 127100 117380
rect 127400 117120 127600 117380
rect 127900 117120 128100 117380
rect 128400 117120 128600 117380
rect 128900 117120 129100 117380
rect 129400 117120 129600 117380
rect 129900 117120 130100 117380
rect 130400 117120 130600 117380
rect 130900 117120 131100 117380
rect 131400 117120 131600 117380
rect 131900 117120 132100 117380
rect 132400 117120 132600 117380
rect 132900 117120 133100 117380
rect 133400 117120 133600 117380
rect 133900 117120 134100 117380
rect 134400 117120 134600 117380
rect 134900 117120 135100 117380
rect 135400 117120 135600 117380
rect 135900 117120 136100 117380
rect 136400 117120 136600 117380
rect 136900 117120 137100 117380
rect 137400 117120 137600 117380
rect 137900 117120 138100 117380
rect 138400 117120 138600 117380
rect 138900 117120 139100 117380
rect 139400 117120 139600 117380
rect 139900 117120 140100 117380
rect 140400 117120 140600 117380
rect 140900 117120 141100 117380
rect 141400 117120 141600 117380
rect 141900 117120 142000 117380
rect 118000 117100 118120 117120
rect 118380 117100 118620 117120
rect 118880 117100 119120 117120
rect 119380 117100 119620 117120
rect 119880 117100 120120 117120
rect 120380 117100 120620 117120
rect 120880 117100 121120 117120
rect 121380 117100 121620 117120
rect 121880 117100 122120 117120
rect 122380 117100 122620 117120
rect 122880 117100 123120 117120
rect 123380 117100 123620 117120
rect 123880 117100 124120 117120
rect 124380 117100 124620 117120
rect 124880 117100 125120 117120
rect 125380 117100 125620 117120
rect 125880 117100 126120 117120
rect 126380 117100 126620 117120
rect 126880 117100 127120 117120
rect 127380 117100 127620 117120
rect 127880 117100 128120 117120
rect 128380 117100 128620 117120
rect 128880 117100 129120 117120
rect 129380 117100 129620 117120
rect 129880 117100 130120 117120
rect 130380 117100 130620 117120
rect 130880 117100 131120 117120
rect 131380 117100 131620 117120
rect 131880 117100 132120 117120
rect 132380 117100 132620 117120
rect 132880 117100 133120 117120
rect 133380 117100 133620 117120
rect 133880 117100 134120 117120
rect 134380 117100 134620 117120
rect 134880 117100 135120 117120
rect 135380 117100 135620 117120
rect 135880 117100 136120 117120
rect 136380 117100 136620 117120
rect 136880 117100 137120 117120
rect 137380 117100 137620 117120
rect 137880 117100 138120 117120
rect 138380 117100 138620 117120
rect 138880 117100 139120 117120
rect 139380 117100 139620 117120
rect 139880 117100 140120 117120
rect 140380 117100 140620 117120
rect 140880 117100 141120 117120
rect 141380 117100 141620 117120
rect 141880 117100 142000 117120
rect 118000 116900 142000 117100
rect 118000 116880 118120 116900
rect 118380 116880 118620 116900
rect 118880 116880 119120 116900
rect 119380 116880 119620 116900
rect 119880 116880 120120 116900
rect 120380 116880 120620 116900
rect 120880 116880 121120 116900
rect 121380 116880 121620 116900
rect 121880 116880 122120 116900
rect 122380 116880 122620 116900
rect 122880 116880 123120 116900
rect 123380 116880 123620 116900
rect 123880 116880 124120 116900
rect 124380 116880 124620 116900
rect 124880 116880 125120 116900
rect 125380 116880 125620 116900
rect 125880 116880 126120 116900
rect 126380 116880 126620 116900
rect 126880 116880 127120 116900
rect 127380 116880 127620 116900
rect 127880 116880 128120 116900
rect 128380 116880 128620 116900
rect 128880 116880 129120 116900
rect 129380 116880 129620 116900
rect 129880 116880 130120 116900
rect 130380 116880 130620 116900
rect 130880 116880 131120 116900
rect 131380 116880 131620 116900
rect 131880 116880 132120 116900
rect 132380 116880 132620 116900
rect 132880 116880 133120 116900
rect 133380 116880 133620 116900
rect 133880 116880 134120 116900
rect 134380 116880 134620 116900
rect 134880 116880 135120 116900
rect 135380 116880 135620 116900
rect 135880 116880 136120 116900
rect 136380 116880 136620 116900
rect 136880 116880 137120 116900
rect 137380 116880 137620 116900
rect 137880 116880 138120 116900
rect 138380 116880 138620 116900
rect 138880 116880 139120 116900
rect 139380 116880 139620 116900
rect 139880 116880 140120 116900
rect 140380 116880 140620 116900
rect 140880 116880 141120 116900
rect 141380 116880 141620 116900
rect 141880 116880 142000 116900
rect 118000 116620 118100 116880
rect 118400 116620 118600 116880
rect 118900 116620 119100 116880
rect 119400 116620 119600 116880
rect 119900 116620 120100 116880
rect 120400 116620 120600 116880
rect 120900 116620 121100 116880
rect 121400 116620 121600 116880
rect 121900 116620 122100 116880
rect 122400 116620 122600 116880
rect 122900 116620 123100 116880
rect 123400 116620 123600 116880
rect 123900 116620 124100 116880
rect 124400 116620 124600 116880
rect 124900 116620 125100 116880
rect 125400 116620 125600 116880
rect 125900 116620 126100 116880
rect 126400 116620 126600 116880
rect 126900 116620 127100 116880
rect 127400 116620 127600 116880
rect 127900 116620 128100 116880
rect 128400 116620 128600 116880
rect 128900 116620 129100 116880
rect 129400 116620 129600 116880
rect 129900 116620 130100 116880
rect 130400 116620 130600 116880
rect 130900 116620 131100 116880
rect 131400 116620 131600 116880
rect 131900 116620 132100 116880
rect 132400 116620 132600 116880
rect 132900 116620 133100 116880
rect 133400 116620 133600 116880
rect 133900 116620 134100 116880
rect 134400 116620 134600 116880
rect 134900 116620 135100 116880
rect 135400 116620 135600 116880
rect 135900 116620 136100 116880
rect 136400 116620 136600 116880
rect 136900 116620 137100 116880
rect 137400 116620 137600 116880
rect 137900 116620 138100 116880
rect 138400 116620 138600 116880
rect 138900 116620 139100 116880
rect 139400 116620 139600 116880
rect 139900 116620 140100 116880
rect 140400 116620 140600 116880
rect 140900 116620 141100 116880
rect 141400 116620 141600 116880
rect 141900 116620 142000 116880
rect 118000 116600 118120 116620
rect 118380 116600 118620 116620
rect 118880 116600 119120 116620
rect 119380 116600 119620 116620
rect 119880 116600 120120 116620
rect 120380 116600 120620 116620
rect 120880 116600 121120 116620
rect 121380 116600 121620 116620
rect 121880 116600 122120 116620
rect 122380 116600 122620 116620
rect 122880 116600 123120 116620
rect 123380 116600 123620 116620
rect 123880 116600 124120 116620
rect 124380 116600 124620 116620
rect 124880 116600 125120 116620
rect 125380 116600 125620 116620
rect 125880 116600 126120 116620
rect 126380 116600 126620 116620
rect 126880 116600 127120 116620
rect 127380 116600 127620 116620
rect 127880 116600 128120 116620
rect 128380 116600 128620 116620
rect 128880 116600 129120 116620
rect 129380 116600 129620 116620
rect 129880 116600 130120 116620
rect 130380 116600 130620 116620
rect 130880 116600 131120 116620
rect 131380 116600 131620 116620
rect 131880 116600 132120 116620
rect 132380 116600 132620 116620
rect 132880 116600 133120 116620
rect 133380 116600 133620 116620
rect 133880 116600 134120 116620
rect 134380 116600 134620 116620
rect 134880 116600 135120 116620
rect 135380 116600 135620 116620
rect 135880 116600 136120 116620
rect 136380 116600 136620 116620
rect 136880 116600 137120 116620
rect 137380 116600 137620 116620
rect 137880 116600 138120 116620
rect 138380 116600 138620 116620
rect 138880 116600 139120 116620
rect 139380 116600 139620 116620
rect 139880 116600 140120 116620
rect 140380 116600 140620 116620
rect 140880 116600 141120 116620
rect 141380 116600 141620 116620
rect 141880 116600 142000 116620
rect 118000 116400 142000 116600
rect 118000 116380 118120 116400
rect 118380 116380 118620 116400
rect 118880 116380 119120 116400
rect 119380 116380 119620 116400
rect 119880 116380 120120 116400
rect 120380 116380 120620 116400
rect 120880 116380 121120 116400
rect 121380 116380 121620 116400
rect 121880 116380 122120 116400
rect 122380 116380 122620 116400
rect 122880 116380 123120 116400
rect 123380 116380 123620 116400
rect 123880 116380 124120 116400
rect 124380 116380 124620 116400
rect 124880 116380 125120 116400
rect 125380 116380 125620 116400
rect 125880 116380 126120 116400
rect 126380 116380 126620 116400
rect 126880 116380 127120 116400
rect 127380 116380 127620 116400
rect 127880 116380 128120 116400
rect 128380 116380 128620 116400
rect 128880 116380 129120 116400
rect 129380 116380 129620 116400
rect 129880 116380 130120 116400
rect 130380 116380 130620 116400
rect 130880 116380 131120 116400
rect 131380 116380 131620 116400
rect 131880 116380 132120 116400
rect 132380 116380 132620 116400
rect 132880 116380 133120 116400
rect 133380 116380 133620 116400
rect 133880 116380 134120 116400
rect 134380 116380 134620 116400
rect 134880 116380 135120 116400
rect 135380 116380 135620 116400
rect 135880 116380 136120 116400
rect 136380 116380 136620 116400
rect 136880 116380 137120 116400
rect 137380 116380 137620 116400
rect 137880 116380 138120 116400
rect 138380 116380 138620 116400
rect 138880 116380 139120 116400
rect 139380 116380 139620 116400
rect 139880 116380 140120 116400
rect 140380 116380 140620 116400
rect 140880 116380 141120 116400
rect 141380 116380 141620 116400
rect 141880 116380 142000 116400
rect 118000 116120 118100 116380
rect 118400 116120 118600 116380
rect 118900 116120 119100 116380
rect 119400 116120 119600 116380
rect 119900 116120 120100 116380
rect 120400 116120 120600 116380
rect 120900 116120 121100 116380
rect 121400 116120 121600 116380
rect 121900 116120 122100 116380
rect 122400 116120 122600 116380
rect 122900 116120 123100 116380
rect 123400 116120 123600 116380
rect 123900 116120 124100 116380
rect 124400 116120 124600 116380
rect 124900 116120 125100 116380
rect 125400 116120 125600 116380
rect 125900 116120 126100 116380
rect 126400 116120 126600 116380
rect 126900 116120 127100 116380
rect 127400 116120 127600 116380
rect 127900 116120 128100 116380
rect 128400 116120 128600 116380
rect 128900 116120 129100 116380
rect 129400 116120 129600 116380
rect 129900 116120 130100 116380
rect 130400 116120 130600 116380
rect 130900 116120 131100 116380
rect 131400 116120 131600 116380
rect 131900 116120 132100 116380
rect 132400 116120 132600 116380
rect 132900 116120 133100 116380
rect 133400 116120 133600 116380
rect 133900 116120 134100 116380
rect 134400 116120 134600 116380
rect 134900 116120 135100 116380
rect 135400 116120 135600 116380
rect 135900 116120 136100 116380
rect 136400 116120 136600 116380
rect 136900 116120 137100 116380
rect 137400 116120 137600 116380
rect 137900 116120 138100 116380
rect 138400 116120 138600 116380
rect 138900 116120 139100 116380
rect 139400 116120 139600 116380
rect 139900 116120 140100 116380
rect 140400 116120 140600 116380
rect 140900 116120 141100 116380
rect 141400 116120 141600 116380
rect 141900 116120 142000 116380
rect 118000 116100 118120 116120
rect 118380 116100 118620 116120
rect 118880 116100 119120 116120
rect 119380 116100 119620 116120
rect 119880 116100 120120 116120
rect 120380 116100 120620 116120
rect 120880 116100 121120 116120
rect 121380 116100 121620 116120
rect 121880 116100 122120 116120
rect 122380 116100 122620 116120
rect 122880 116100 123120 116120
rect 123380 116100 123620 116120
rect 123880 116100 124120 116120
rect 124380 116100 124620 116120
rect 124880 116100 125120 116120
rect 125380 116100 125620 116120
rect 125880 116100 126120 116120
rect 126380 116100 126620 116120
rect 126880 116100 127120 116120
rect 127380 116100 127620 116120
rect 127880 116100 128120 116120
rect 128380 116100 128620 116120
rect 128880 116100 129120 116120
rect 129380 116100 129620 116120
rect 129880 116100 130120 116120
rect 130380 116100 130620 116120
rect 130880 116100 131120 116120
rect 131380 116100 131620 116120
rect 131880 116100 132120 116120
rect 132380 116100 132620 116120
rect 132880 116100 133120 116120
rect 133380 116100 133620 116120
rect 133880 116100 134120 116120
rect 134380 116100 134620 116120
rect 134880 116100 135120 116120
rect 135380 116100 135620 116120
rect 135880 116100 136120 116120
rect 136380 116100 136620 116120
rect 136880 116100 137120 116120
rect 137380 116100 137620 116120
rect 137880 116100 138120 116120
rect 138380 116100 138620 116120
rect 138880 116100 139120 116120
rect 139380 116100 139620 116120
rect 139880 116100 140120 116120
rect 140380 116100 140620 116120
rect 140880 116100 141120 116120
rect 141380 116100 141620 116120
rect 141880 116100 142000 116120
rect 118000 115900 142000 116100
rect 118000 115880 118120 115900
rect 118380 115880 118620 115900
rect 118880 115880 119120 115900
rect 119380 115880 119620 115900
rect 119880 115880 120120 115900
rect 120380 115880 120620 115900
rect 120880 115880 121120 115900
rect 121380 115880 121620 115900
rect 121880 115880 122120 115900
rect 122380 115880 122620 115900
rect 122880 115880 123120 115900
rect 123380 115880 123620 115900
rect 123880 115880 124120 115900
rect 124380 115880 124620 115900
rect 124880 115880 125120 115900
rect 125380 115880 125620 115900
rect 125880 115880 126120 115900
rect 126380 115880 126620 115900
rect 126880 115880 127120 115900
rect 127380 115880 127620 115900
rect 127880 115880 128120 115900
rect 128380 115880 128620 115900
rect 128880 115880 129120 115900
rect 129380 115880 129620 115900
rect 129880 115880 130120 115900
rect 130380 115880 130620 115900
rect 130880 115880 131120 115900
rect 131380 115880 131620 115900
rect 131880 115880 132120 115900
rect 132380 115880 132620 115900
rect 132880 115880 133120 115900
rect 133380 115880 133620 115900
rect 133880 115880 134120 115900
rect 134380 115880 134620 115900
rect 134880 115880 135120 115900
rect 135380 115880 135620 115900
rect 135880 115880 136120 115900
rect 136380 115880 136620 115900
rect 136880 115880 137120 115900
rect 137380 115880 137620 115900
rect 137880 115880 138120 115900
rect 138380 115880 138620 115900
rect 138880 115880 139120 115900
rect 139380 115880 139620 115900
rect 139880 115880 140120 115900
rect 140380 115880 140620 115900
rect 140880 115880 141120 115900
rect 141380 115880 141620 115900
rect 141880 115880 142000 115900
rect 118000 115620 118100 115880
rect 118400 115620 118600 115880
rect 118900 115620 119100 115880
rect 119400 115620 119600 115880
rect 119900 115620 120100 115880
rect 120400 115620 120600 115880
rect 120900 115620 121100 115880
rect 121400 115620 121600 115880
rect 121900 115620 122100 115880
rect 122400 115620 122600 115880
rect 122900 115620 123100 115880
rect 123400 115620 123600 115880
rect 123900 115620 124100 115880
rect 124400 115620 124600 115880
rect 124900 115620 125100 115880
rect 125400 115620 125600 115880
rect 125900 115620 126100 115880
rect 126400 115620 126600 115880
rect 126900 115620 127100 115880
rect 127400 115620 127600 115880
rect 127900 115620 128100 115880
rect 128400 115620 128600 115880
rect 128900 115620 129100 115880
rect 129400 115620 129600 115880
rect 129900 115620 130100 115880
rect 130400 115620 130600 115880
rect 130900 115620 131100 115880
rect 131400 115620 131600 115880
rect 131900 115620 132100 115880
rect 132400 115620 132600 115880
rect 132900 115620 133100 115880
rect 133400 115620 133600 115880
rect 133900 115620 134100 115880
rect 134400 115620 134600 115880
rect 134900 115620 135100 115880
rect 135400 115620 135600 115880
rect 135900 115620 136100 115880
rect 136400 115620 136600 115880
rect 136900 115620 137100 115880
rect 137400 115620 137600 115880
rect 137900 115620 138100 115880
rect 138400 115620 138600 115880
rect 138900 115620 139100 115880
rect 139400 115620 139600 115880
rect 139900 115620 140100 115880
rect 140400 115620 140600 115880
rect 140900 115620 141100 115880
rect 141400 115620 141600 115880
rect 141900 115620 142000 115880
rect 118000 115600 118120 115620
rect 118380 115600 118620 115620
rect 118880 115600 119120 115620
rect 119380 115600 119620 115620
rect 119880 115600 120120 115620
rect 120380 115600 120620 115620
rect 120880 115600 121120 115620
rect 121380 115600 121620 115620
rect 121880 115600 122120 115620
rect 122380 115600 122620 115620
rect 122880 115600 123120 115620
rect 123380 115600 123620 115620
rect 123880 115600 124120 115620
rect 124380 115600 124620 115620
rect 124880 115600 125120 115620
rect 125380 115600 125620 115620
rect 125880 115600 126120 115620
rect 126380 115600 126620 115620
rect 126880 115600 127120 115620
rect 127380 115600 127620 115620
rect 127880 115600 128120 115620
rect 128380 115600 128620 115620
rect 128880 115600 129120 115620
rect 129380 115600 129620 115620
rect 129880 115600 130120 115620
rect 130380 115600 130620 115620
rect 130880 115600 131120 115620
rect 131380 115600 131620 115620
rect 131880 115600 132120 115620
rect 132380 115600 132620 115620
rect 132880 115600 133120 115620
rect 133380 115600 133620 115620
rect 133880 115600 134120 115620
rect 134380 115600 134620 115620
rect 134880 115600 135120 115620
rect 135380 115600 135620 115620
rect 135880 115600 136120 115620
rect 136380 115600 136620 115620
rect 136880 115600 137120 115620
rect 137380 115600 137620 115620
rect 137880 115600 138120 115620
rect 138380 115600 138620 115620
rect 138880 115600 139120 115620
rect 139380 115600 139620 115620
rect 139880 115600 140120 115620
rect 140380 115600 140620 115620
rect 140880 115600 141120 115620
rect 141380 115600 141620 115620
rect 141880 115600 142000 115620
rect 118000 115400 142000 115600
rect 118000 115380 118120 115400
rect 118380 115380 118620 115400
rect 118880 115380 119120 115400
rect 119380 115380 119620 115400
rect 119880 115380 120120 115400
rect 120380 115380 120620 115400
rect 120880 115380 121120 115400
rect 121380 115380 121620 115400
rect 121880 115380 122120 115400
rect 122380 115380 122620 115400
rect 122880 115380 123120 115400
rect 123380 115380 123620 115400
rect 123880 115380 124120 115400
rect 124380 115380 124620 115400
rect 124880 115380 125120 115400
rect 125380 115380 125620 115400
rect 125880 115380 126120 115400
rect 126380 115380 126620 115400
rect 126880 115380 127120 115400
rect 127380 115380 127620 115400
rect 127880 115380 128120 115400
rect 128380 115380 128620 115400
rect 128880 115380 129120 115400
rect 129380 115380 129620 115400
rect 129880 115380 130120 115400
rect 130380 115380 130620 115400
rect 130880 115380 131120 115400
rect 131380 115380 131620 115400
rect 131880 115380 132120 115400
rect 132380 115380 132620 115400
rect 132880 115380 133120 115400
rect 133380 115380 133620 115400
rect 133880 115380 134120 115400
rect 134380 115380 134620 115400
rect 134880 115380 135120 115400
rect 135380 115380 135620 115400
rect 135880 115380 136120 115400
rect 136380 115380 136620 115400
rect 136880 115380 137120 115400
rect 137380 115380 137620 115400
rect 137880 115380 138120 115400
rect 138380 115380 138620 115400
rect 138880 115380 139120 115400
rect 139380 115380 139620 115400
rect 139880 115380 140120 115400
rect 140380 115380 140620 115400
rect 140880 115380 141120 115400
rect 141380 115380 141620 115400
rect 141880 115380 142000 115400
rect 118000 115120 118100 115380
rect 118400 115120 118600 115380
rect 118900 115120 119100 115380
rect 119400 115120 119600 115380
rect 119900 115120 120100 115380
rect 120400 115120 120600 115380
rect 120900 115120 121100 115380
rect 121400 115120 121600 115380
rect 121900 115120 122100 115380
rect 122400 115120 122600 115380
rect 122900 115120 123100 115380
rect 123400 115120 123600 115380
rect 123900 115120 124100 115380
rect 124400 115120 124600 115380
rect 124900 115120 125100 115380
rect 125400 115120 125600 115380
rect 125900 115120 126100 115380
rect 126400 115120 126600 115380
rect 126900 115120 127100 115380
rect 127400 115120 127600 115380
rect 127900 115120 128100 115380
rect 128400 115120 128600 115380
rect 128900 115120 129100 115380
rect 129400 115120 129600 115380
rect 129900 115120 130100 115380
rect 130400 115120 130600 115380
rect 130900 115120 131100 115380
rect 131400 115120 131600 115380
rect 131900 115120 132100 115380
rect 132400 115120 132600 115380
rect 132900 115120 133100 115380
rect 133400 115120 133600 115380
rect 133900 115120 134100 115380
rect 134400 115120 134600 115380
rect 134900 115120 135100 115380
rect 135400 115120 135600 115380
rect 135900 115120 136100 115380
rect 136400 115120 136600 115380
rect 136900 115120 137100 115380
rect 137400 115120 137600 115380
rect 137900 115120 138100 115380
rect 138400 115120 138600 115380
rect 138900 115120 139100 115380
rect 139400 115120 139600 115380
rect 139900 115120 140100 115380
rect 140400 115120 140600 115380
rect 140900 115120 141100 115380
rect 141400 115120 141600 115380
rect 141900 115120 142000 115380
rect 118000 115100 118120 115120
rect 118380 115100 118620 115120
rect 118880 115100 119120 115120
rect 119380 115100 119620 115120
rect 119880 115100 120120 115120
rect 120380 115100 120620 115120
rect 120880 115100 121120 115120
rect 121380 115100 121620 115120
rect 121880 115100 122120 115120
rect 122380 115100 122620 115120
rect 122880 115100 123120 115120
rect 123380 115100 123620 115120
rect 123880 115100 124120 115120
rect 124380 115100 124620 115120
rect 124880 115100 125120 115120
rect 125380 115100 125620 115120
rect 125880 115100 126120 115120
rect 126380 115100 126620 115120
rect 126880 115100 127120 115120
rect 127380 115100 127620 115120
rect 127880 115100 128120 115120
rect 128380 115100 128620 115120
rect 128880 115100 129120 115120
rect 129380 115100 129620 115120
rect 129880 115100 130120 115120
rect 130380 115100 130620 115120
rect 130880 115100 131120 115120
rect 131380 115100 131620 115120
rect 131880 115100 132120 115120
rect 132380 115100 132620 115120
rect 132880 115100 133120 115120
rect 133380 115100 133620 115120
rect 133880 115100 134120 115120
rect 134380 115100 134620 115120
rect 134880 115100 135120 115120
rect 135380 115100 135620 115120
rect 135880 115100 136120 115120
rect 136380 115100 136620 115120
rect 136880 115100 137120 115120
rect 137380 115100 137620 115120
rect 137880 115100 138120 115120
rect 138380 115100 138620 115120
rect 138880 115100 139120 115120
rect 139380 115100 139620 115120
rect 139880 115100 140120 115120
rect 140380 115100 140620 115120
rect 140880 115100 141120 115120
rect 141380 115100 141620 115120
rect 141880 115100 142000 115120
rect 118000 114900 142000 115100
rect 118000 114880 118120 114900
rect 118380 114880 118620 114900
rect 118880 114880 119120 114900
rect 119380 114880 119620 114900
rect 119880 114880 120120 114900
rect 120380 114880 120620 114900
rect 120880 114880 121120 114900
rect 121380 114880 121620 114900
rect 121880 114880 122120 114900
rect 122380 114880 122620 114900
rect 122880 114880 123120 114900
rect 123380 114880 123620 114900
rect 123880 114880 124120 114900
rect 124380 114880 124620 114900
rect 124880 114880 125120 114900
rect 125380 114880 125620 114900
rect 125880 114880 126120 114900
rect 126380 114880 126620 114900
rect 126880 114880 127120 114900
rect 127380 114880 127620 114900
rect 127880 114880 128120 114900
rect 128380 114880 128620 114900
rect 128880 114880 129120 114900
rect 129380 114880 129620 114900
rect 129880 114880 130120 114900
rect 130380 114880 130620 114900
rect 130880 114880 131120 114900
rect 131380 114880 131620 114900
rect 131880 114880 132120 114900
rect 132380 114880 132620 114900
rect 132880 114880 133120 114900
rect 133380 114880 133620 114900
rect 133880 114880 134120 114900
rect 134380 114880 134620 114900
rect 134880 114880 135120 114900
rect 135380 114880 135620 114900
rect 135880 114880 136120 114900
rect 136380 114880 136620 114900
rect 136880 114880 137120 114900
rect 137380 114880 137620 114900
rect 137880 114880 138120 114900
rect 138380 114880 138620 114900
rect 138880 114880 139120 114900
rect 139380 114880 139620 114900
rect 139880 114880 140120 114900
rect 140380 114880 140620 114900
rect 140880 114880 141120 114900
rect 141380 114880 141620 114900
rect 141880 114880 142000 114900
rect 118000 114620 118100 114880
rect 118400 114620 118600 114880
rect 118900 114620 119100 114880
rect 119400 114620 119600 114880
rect 119900 114620 120100 114880
rect 120400 114620 120600 114880
rect 120900 114620 121100 114880
rect 121400 114620 121600 114880
rect 121900 114620 122100 114880
rect 122400 114620 122600 114880
rect 122900 114620 123100 114880
rect 123400 114620 123600 114880
rect 123900 114620 124100 114880
rect 124400 114620 124600 114880
rect 124900 114620 125100 114880
rect 125400 114620 125600 114880
rect 125900 114620 126100 114880
rect 126400 114620 126600 114880
rect 126900 114620 127100 114880
rect 127400 114620 127600 114880
rect 127900 114620 128100 114880
rect 128400 114620 128600 114880
rect 128900 114620 129100 114880
rect 129400 114620 129600 114880
rect 129900 114620 130100 114880
rect 130400 114620 130600 114880
rect 130900 114620 131100 114880
rect 131400 114620 131600 114880
rect 131900 114620 132100 114880
rect 132400 114620 132600 114880
rect 132900 114620 133100 114880
rect 133400 114620 133600 114880
rect 133900 114620 134100 114880
rect 134400 114620 134600 114880
rect 134900 114620 135100 114880
rect 135400 114620 135600 114880
rect 135900 114620 136100 114880
rect 136400 114620 136600 114880
rect 136900 114620 137100 114880
rect 137400 114620 137600 114880
rect 137900 114620 138100 114880
rect 138400 114620 138600 114880
rect 138900 114620 139100 114880
rect 139400 114620 139600 114880
rect 139900 114620 140100 114880
rect 140400 114620 140600 114880
rect 140900 114620 141100 114880
rect 141400 114620 141600 114880
rect 141900 114620 142000 114880
rect 118000 114600 118120 114620
rect 118380 114600 118620 114620
rect 118880 114600 119120 114620
rect 119380 114600 119620 114620
rect 119880 114600 120120 114620
rect 120380 114600 120620 114620
rect 120880 114600 121120 114620
rect 121380 114600 121620 114620
rect 121880 114600 122120 114620
rect 122380 114600 122620 114620
rect 122880 114600 123120 114620
rect 123380 114600 123620 114620
rect 123880 114600 124120 114620
rect 124380 114600 124620 114620
rect 124880 114600 125120 114620
rect 125380 114600 125620 114620
rect 125880 114600 126120 114620
rect 126380 114600 126620 114620
rect 126880 114600 127120 114620
rect 127380 114600 127620 114620
rect 127880 114600 128120 114620
rect 128380 114600 128620 114620
rect 128880 114600 129120 114620
rect 129380 114600 129620 114620
rect 129880 114600 130120 114620
rect 130380 114600 130620 114620
rect 130880 114600 131120 114620
rect 131380 114600 131620 114620
rect 131880 114600 132120 114620
rect 132380 114600 132620 114620
rect 132880 114600 133120 114620
rect 133380 114600 133620 114620
rect 133880 114600 134120 114620
rect 134380 114600 134620 114620
rect 134880 114600 135120 114620
rect 135380 114600 135620 114620
rect 135880 114600 136120 114620
rect 136380 114600 136620 114620
rect 136880 114600 137120 114620
rect 137380 114600 137620 114620
rect 137880 114600 138120 114620
rect 138380 114600 138620 114620
rect 138880 114600 139120 114620
rect 139380 114600 139620 114620
rect 139880 114600 140120 114620
rect 140380 114600 140620 114620
rect 140880 114600 141120 114620
rect 141380 114600 141620 114620
rect 141880 114600 142000 114620
rect 118000 114400 142000 114600
rect 118000 114380 118120 114400
rect 118380 114380 118620 114400
rect 118880 114380 119120 114400
rect 119380 114380 119620 114400
rect 119880 114380 120120 114400
rect 120380 114380 120620 114400
rect 120880 114380 121120 114400
rect 121380 114380 121620 114400
rect 121880 114380 122120 114400
rect 122380 114380 122620 114400
rect 122880 114380 123120 114400
rect 123380 114380 123620 114400
rect 123880 114380 124120 114400
rect 124380 114380 124620 114400
rect 124880 114380 125120 114400
rect 125380 114380 125620 114400
rect 125880 114380 126120 114400
rect 126380 114380 126620 114400
rect 126880 114380 127120 114400
rect 127380 114380 127620 114400
rect 127880 114380 128120 114400
rect 128380 114380 128620 114400
rect 128880 114380 129120 114400
rect 129380 114380 129620 114400
rect 129880 114380 130120 114400
rect 130380 114380 130620 114400
rect 130880 114380 131120 114400
rect 131380 114380 131620 114400
rect 131880 114380 132120 114400
rect 132380 114380 132620 114400
rect 132880 114380 133120 114400
rect 133380 114380 133620 114400
rect 133880 114380 134120 114400
rect 134380 114380 134620 114400
rect 134880 114380 135120 114400
rect 135380 114380 135620 114400
rect 135880 114380 136120 114400
rect 136380 114380 136620 114400
rect 136880 114380 137120 114400
rect 137380 114380 137620 114400
rect 137880 114380 138120 114400
rect 138380 114380 138620 114400
rect 138880 114380 139120 114400
rect 139380 114380 139620 114400
rect 139880 114380 140120 114400
rect 140380 114380 140620 114400
rect 140880 114380 141120 114400
rect 141380 114380 141620 114400
rect 141880 114380 142000 114400
rect 118000 114120 118100 114380
rect 118400 114120 118600 114380
rect 118900 114120 119100 114380
rect 119400 114120 119600 114380
rect 119900 114120 120100 114380
rect 120400 114120 120600 114380
rect 120900 114120 121100 114380
rect 121400 114120 121600 114380
rect 121900 114120 122100 114380
rect 122400 114120 122600 114380
rect 122900 114120 123100 114380
rect 123400 114120 123600 114380
rect 123900 114120 124100 114380
rect 124400 114120 124600 114380
rect 124900 114120 125100 114380
rect 125400 114120 125600 114380
rect 125900 114120 126100 114380
rect 126400 114120 126600 114380
rect 126900 114120 127100 114380
rect 127400 114120 127600 114380
rect 127900 114120 128100 114380
rect 128400 114120 128600 114380
rect 128900 114120 129100 114380
rect 129400 114120 129600 114380
rect 129900 114120 130100 114380
rect 130400 114120 130600 114380
rect 130900 114120 131100 114380
rect 131400 114120 131600 114380
rect 131900 114120 132100 114380
rect 132400 114120 132600 114380
rect 132900 114120 133100 114380
rect 133400 114120 133600 114380
rect 133900 114120 134100 114380
rect 134400 114120 134600 114380
rect 134900 114120 135100 114380
rect 135400 114120 135600 114380
rect 135900 114120 136100 114380
rect 136400 114120 136600 114380
rect 136900 114120 137100 114380
rect 137400 114120 137600 114380
rect 137900 114120 138100 114380
rect 138400 114120 138600 114380
rect 138900 114120 139100 114380
rect 139400 114120 139600 114380
rect 139900 114120 140100 114380
rect 140400 114120 140600 114380
rect 140900 114120 141100 114380
rect 141400 114120 141600 114380
rect 141900 114120 142000 114380
rect 118000 114100 118120 114120
rect 118380 114100 118620 114120
rect 118880 114100 119120 114120
rect 119380 114100 119620 114120
rect 119880 114100 120120 114120
rect 120380 114100 120620 114120
rect 120880 114100 121120 114120
rect 121380 114100 121620 114120
rect 121880 114100 122120 114120
rect 122380 114100 122620 114120
rect 122880 114100 123120 114120
rect 123380 114100 123620 114120
rect 123880 114100 124120 114120
rect 124380 114100 124620 114120
rect 124880 114100 125120 114120
rect 125380 114100 125620 114120
rect 125880 114100 126120 114120
rect 126380 114100 126620 114120
rect 126880 114100 127120 114120
rect 127380 114100 127620 114120
rect 127880 114100 128120 114120
rect 128380 114100 128620 114120
rect 128880 114100 129120 114120
rect 129380 114100 129620 114120
rect 129880 114100 130120 114120
rect 130380 114100 130620 114120
rect 130880 114100 131120 114120
rect 131380 114100 131620 114120
rect 131880 114100 132120 114120
rect 132380 114100 132620 114120
rect 132880 114100 133120 114120
rect 133380 114100 133620 114120
rect 133880 114100 134120 114120
rect 134380 114100 134620 114120
rect 134880 114100 135120 114120
rect 135380 114100 135620 114120
rect 135880 114100 136120 114120
rect 136380 114100 136620 114120
rect 136880 114100 137120 114120
rect 137380 114100 137620 114120
rect 137880 114100 138120 114120
rect 138380 114100 138620 114120
rect 138880 114100 139120 114120
rect 139380 114100 139620 114120
rect 139880 114100 140120 114120
rect 140380 114100 140620 114120
rect 140880 114100 141120 114120
rect 141380 114100 141620 114120
rect 141880 114100 142000 114120
rect 118000 114000 142000 114100
rect 162000 121900 184000 122000
rect 162000 121880 162120 121900
rect 162380 121880 162620 121900
rect 162880 121880 163120 121900
rect 163380 121880 163620 121900
rect 163880 121880 164120 121900
rect 164380 121880 164620 121900
rect 164880 121880 165120 121900
rect 165380 121880 165620 121900
rect 165880 121880 166120 121900
rect 166380 121880 166620 121900
rect 166880 121880 167120 121900
rect 167380 121880 167620 121900
rect 167880 121880 168120 121900
rect 168380 121880 168620 121900
rect 168880 121880 169120 121900
rect 169380 121880 169620 121900
rect 169880 121880 170120 121900
rect 170380 121880 170620 121900
rect 170880 121880 182120 121900
rect 182380 121880 182620 121900
rect 182880 121880 183120 121900
rect 183380 121880 183620 121900
rect 183880 121880 184000 121900
rect 162000 121620 162100 121880
rect 162400 121620 162600 121880
rect 162900 121620 163100 121880
rect 163400 121620 163600 121880
rect 163900 121620 164100 121880
rect 164400 121620 164600 121880
rect 164900 121620 165100 121880
rect 165400 121620 165600 121880
rect 165900 121620 166100 121880
rect 166400 121620 166600 121880
rect 166900 121620 167100 121880
rect 167400 121620 167600 121880
rect 167900 121620 168100 121880
rect 168400 121620 168600 121880
rect 168900 121620 169100 121880
rect 169400 121620 169600 121880
rect 169900 121620 170100 121880
rect 170400 121620 170600 121880
rect 170900 121800 182100 121880
rect 170900 121620 171200 121800
rect 162000 121600 162120 121620
rect 162380 121600 162620 121620
rect 162880 121600 163120 121620
rect 163380 121600 163620 121620
rect 163880 121600 164120 121620
rect 164380 121600 164620 121620
rect 164880 121600 165120 121620
rect 165380 121600 165620 121620
rect 165880 121600 166120 121620
rect 166380 121600 166620 121620
rect 166880 121600 167120 121620
rect 167380 121600 167620 121620
rect 167880 121600 168120 121620
rect 168380 121600 168620 121620
rect 168880 121600 169120 121620
rect 169380 121600 169620 121620
rect 169880 121600 170120 121620
rect 170380 121600 170620 121620
rect 170880 121600 171200 121620
rect 162000 121400 171200 121600
rect 162000 121380 162120 121400
rect 162380 121380 162620 121400
rect 162880 121380 163120 121400
rect 163380 121380 163620 121400
rect 163880 121380 164120 121400
rect 164380 121380 164620 121400
rect 164880 121380 165120 121400
rect 165380 121380 165620 121400
rect 165880 121380 166120 121400
rect 166380 121380 166620 121400
rect 166880 121380 167120 121400
rect 167380 121380 167620 121400
rect 167880 121380 168120 121400
rect 168380 121380 168620 121400
rect 168880 121380 169120 121400
rect 169380 121380 169620 121400
rect 169880 121380 170120 121400
rect 170380 121380 170620 121400
rect 170880 121380 171200 121400
rect 162000 121120 162100 121380
rect 162400 121120 162600 121380
rect 162900 121120 163100 121380
rect 163400 121120 163600 121380
rect 163900 121120 164100 121380
rect 164400 121120 164600 121380
rect 164900 121120 165100 121380
rect 165400 121120 165600 121380
rect 165900 121120 166100 121380
rect 166400 121120 166600 121380
rect 166900 121120 167100 121380
rect 167400 121120 167600 121380
rect 167900 121120 168100 121380
rect 168400 121120 168600 121380
rect 168900 121120 169100 121380
rect 169400 121120 169600 121380
rect 169900 121120 170100 121380
rect 170400 121120 170600 121380
rect 170900 121120 171200 121380
rect 162000 121100 162120 121120
rect 162380 121100 162620 121120
rect 162880 121100 163120 121120
rect 163380 121100 163620 121120
rect 163880 121100 164120 121120
rect 164380 121100 164620 121120
rect 164880 121100 165120 121120
rect 165380 121100 165620 121120
rect 165880 121100 166120 121120
rect 166380 121100 166620 121120
rect 166880 121100 167120 121120
rect 167380 121100 167620 121120
rect 167880 121100 168120 121120
rect 168380 121100 168620 121120
rect 168880 121100 169120 121120
rect 169380 121100 169620 121120
rect 169880 121100 170120 121120
rect 170380 121100 170620 121120
rect 170880 121100 171200 121120
rect 162000 120900 171200 121100
rect 162000 120880 162120 120900
rect 162380 120880 162620 120900
rect 162880 120880 163120 120900
rect 163380 120880 163620 120900
rect 163880 120880 164120 120900
rect 164380 120880 164620 120900
rect 164880 120880 165120 120900
rect 165380 120880 165620 120900
rect 165880 120880 166120 120900
rect 166380 120880 166620 120900
rect 166880 120880 167120 120900
rect 167380 120880 167620 120900
rect 167880 120880 168120 120900
rect 168380 120880 168620 120900
rect 168880 120880 169120 120900
rect 169380 120880 169620 120900
rect 169880 120880 170120 120900
rect 170380 120880 170620 120900
rect 170880 120880 171200 120900
rect 162000 120620 162100 120880
rect 162400 120620 162600 120880
rect 162900 120620 163100 120880
rect 163400 120620 163600 120880
rect 163900 120620 164100 120880
rect 164400 120620 164600 120880
rect 164900 120620 165100 120880
rect 165400 120620 165600 120880
rect 165900 120620 166100 120880
rect 166400 120620 166600 120880
rect 166900 120620 167100 120880
rect 167400 120620 167600 120880
rect 167900 120620 168100 120880
rect 168400 120620 168600 120880
rect 168900 120620 169100 120880
rect 169400 120620 169600 120880
rect 169900 120620 170100 120880
rect 170400 120620 170600 120880
rect 170900 120620 171200 120880
rect 162000 120600 162120 120620
rect 162380 120600 162620 120620
rect 162880 120600 163120 120620
rect 163380 120600 163620 120620
rect 163880 120600 164120 120620
rect 164380 120600 164620 120620
rect 164880 120600 165120 120620
rect 165380 120600 165620 120620
rect 165880 120600 166120 120620
rect 166380 120600 166620 120620
rect 166880 120600 167120 120620
rect 167380 120600 167620 120620
rect 167880 120600 168120 120620
rect 168380 120600 168620 120620
rect 168880 120600 169120 120620
rect 169380 120600 169620 120620
rect 169880 120600 170120 120620
rect 170380 120600 170620 120620
rect 170880 120600 171200 120620
rect 162000 120400 171200 120600
rect 162000 120380 162120 120400
rect 162380 120380 162620 120400
rect 162880 120380 163120 120400
rect 163380 120380 163620 120400
rect 163880 120380 164120 120400
rect 164380 120380 164620 120400
rect 164880 120380 165120 120400
rect 165380 120380 165620 120400
rect 165880 120380 166120 120400
rect 166380 120380 166620 120400
rect 166880 120380 167120 120400
rect 167380 120380 167620 120400
rect 167880 120380 168120 120400
rect 168380 120380 168620 120400
rect 168880 120380 169120 120400
rect 169380 120380 169620 120400
rect 169880 120380 170120 120400
rect 170380 120380 170620 120400
rect 170880 120380 171200 120400
rect 162000 120120 162100 120380
rect 162400 120120 162600 120380
rect 162900 120120 163100 120380
rect 163400 120120 163600 120380
rect 163900 120120 164100 120380
rect 164400 120120 164600 120380
rect 164900 120120 165100 120380
rect 165400 120120 165600 120380
rect 165900 120120 166100 120380
rect 166400 120120 166600 120380
rect 166900 120120 167100 120380
rect 167400 120120 167600 120380
rect 167900 120120 168100 120380
rect 168400 120120 168600 120380
rect 168900 120120 169100 120380
rect 169400 120120 169600 120380
rect 169900 120120 170100 120380
rect 170400 120120 170600 120380
rect 170900 120120 171200 120380
rect 162000 120100 162120 120120
rect 162380 120100 162620 120120
rect 162880 120100 163120 120120
rect 163380 120100 163620 120120
rect 163880 120100 164120 120120
rect 164380 120100 164620 120120
rect 164880 120100 165120 120120
rect 165380 120100 165620 120120
rect 165880 120100 166120 120120
rect 166380 120100 166620 120120
rect 166880 120100 167120 120120
rect 167380 120100 167620 120120
rect 167880 120100 168120 120120
rect 168380 120100 168620 120120
rect 168880 120100 169120 120120
rect 169380 120100 169620 120120
rect 169880 120100 170120 120120
rect 170380 120100 170620 120120
rect 170880 120100 171200 120120
rect 162000 119900 171200 120100
rect 162000 119880 162120 119900
rect 162380 119880 162620 119900
rect 162880 119880 163120 119900
rect 163380 119880 163620 119900
rect 163880 119880 164120 119900
rect 164380 119880 164620 119900
rect 164880 119880 165120 119900
rect 165380 119880 165620 119900
rect 165880 119880 166120 119900
rect 166380 119880 166620 119900
rect 166880 119880 167120 119900
rect 167380 119880 167620 119900
rect 167880 119880 168120 119900
rect 168380 119880 168620 119900
rect 168880 119880 169120 119900
rect 169380 119880 169620 119900
rect 169880 119880 170120 119900
rect 170380 119880 170620 119900
rect 170880 119880 171200 119900
rect 162000 119620 162100 119880
rect 162400 119620 162600 119880
rect 162900 119620 163100 119880
rect 163400 119620 163600 119880
rect 163900 119620 164100 119880
rect 164400 119620 164600 119880
rect 164900 119620 165100 119880
rect 165400 119620 165600 119880
rect 165900 119620 166100 119880
rect 166400 119620 166600 119880
rect 166900 119620 167100 119880
rect 167400 119620 167600 119880
rect 167900 119620 168100 119880
rect 168400 119620 168600 119880
rect 168900 119620 169100 119880
rect 169400 119620 169600 119880
rect 169900 119620 170100 119880
rect 170400 119620 170600 119880
rect 170900 119620 171200 119880
rect 162000 119600 162120 119620
rect 162380 119600 162620 119620
rect 162880 119600 163120 119620
rect 163380 119600 163620 119620
rect 163880 119600 164120 119620
rect 164380 119600 164620 119620
rect 164880 119600 165120 119620
rect 165380 119600 165620 119620
rect 165880 119600 166120 119620
rect 166380 119600 166620 119620
rect 166880 119600 167120 119620
rect 167380 119600 167620 119620
rect 167880 119600 168120 119620
rect 168380 119600 168620 119620
rect 168880 119600 169120 119620
rect 169380 119600 169620 119620
rect 169880 119600 170120 119620
rect 170380 119600 170620 119620
rect 170880 119600 171200 119620
rect 181800 121620 182100 121800
rect 182400 121620 182600 121880
rect 182900 121620 183100 121880
rect 183400 121620 183600 121880
rect 183900 121620 184000 121880
rect 181800 121600 182120 121620
rect 182380 121600 182620 121620
rect 182880 121600 183120 121620
rect 183380 121600 183620 121620
rect 183880 121600 184000 121620
rect 181800 121400 184000 121600
rect 181800 121380 182120 121400
rect 182380 121380 182620 121400
rect 182880 121380 183120 121400
rect 183380 121380 183620 121400
rect 183880 121380 184000 121400
rect 181800 121120 182100 121380
rect 182400 121120 182600 121380
rect 182900 121120 183100 121380
rect 183400 121120 183600 121380
rect 183900 121120 184000 121380
rect 181800 121100 182120 121120
rect 182380 121100 182620 121120
rect 182880 121100 183120 121120
rect 183380 121100 183620 121120
rect 183880 121100 184000 121120
rect 181800 120900 184000 121100
rect 181800 120880 182120 120900
rect 182380 120880 182620 120900
rect 182880 120880 183120 120900
rect 183380 120880 183620 120900
rect 183880 120880 184000 120900
rect 181800 120620 182100 120880
rect 182400 120620 182600 120880
rect 182900 120620 183100 120880
rect 183400 120620 183600 120880
rect 183900 120620 184000 120880
rect 181800 120600 182120 120620
rect 182380 120600 182620 120620
rect 182880 120600 183120 120620
rect 183380 120600 183620 120620
rect 183880 120600 184000 120620
rect 181800 120400 184000 120600
rect 181800 120380 182120 120400
rect 182380 120380 182620 120400
rect 182880 120380 183120 120400
rect 183380 120380 183620 120400
rect 183880 120380 184000 120400
rect 181800 120120 182100 120380
rect 182400 120120 182600 120380
rect 182900 120120 183100 120380
rect 183400 120120 183600 120380
rect 183900 120120 184000 120380
rect 181800 120100 182120 120120
rect 182380 120100 182620 120120
rect 182880 120100 183120 120120
rect 183380 120100 183620 120120
rect 183880 120100 184000 120120
rect 181800 119900 184000 120100
rect 181800 119880 182120 119900
rect 182380 119880 182620 119900
rect 182880 119880 183120 119900
rect 183380 119880 183620 119900
rect 183880 119880 184000 119900
rect 181800 119620 182100 119880
rect 182400 119620 182600 119880
rect 182900 119620 183100 119880
rect 183400 119620 183600 119880
rect 183900 119620 184000 119880
rect 181800 119600 182120 119620
rect 182380 119600 182620 119620
rect 182880 119600 183120 119620
rect 183380 119600 183620 119620
rect 183880 119600 184000 119620
rect 162000 119400 184000 119600
rect 162000 119380 162120 119400
rect 162380 119380 162620 119400
rect 162880 119380 163120 119400
rect 163380 119380 163620 119400
rect 163880 119380 164120 119400
rect 164380 119380 164620 119400
rect 164880 119380 165120 119400
rect 165380 119380 165620 119400
rect 165880 119380 166120 119400
rect 166380 119380 166620 119400
rect 166880 119380 167120 119400
rect 167380 119380 167620 119400
rect 167880 119380 168120 119400
rect 168380 119380 168620 119400
rect 168880 119380 169120 119400
rect 169380 119380 169620 119400
rect 169880 119380 170120 119400
rect 170380 119380 170620 119400
rect 170880 119380 171120 119400
rect 171380 119380 171620 119400
rect 171880 119380 172120 119400
rect 172380 119380 172620 119400
rect 172880 119380 173120 119400
rect 173380 119380 173620 119400
rect 173880 119380 174120 119400
rect 174380 119380 174620 119400
rect 174880 119380 175120 119400
rect 175380 119380 175620 119400
rect 175880 119380 176120 119400
rect 176380 119380 176620 119400
rect 176880 119380 177120 119400
rect 177380 119380 177620 119400
rect 177880 119380 178120 119400
rect 178380 119380 178620 119400
rect 178880 119380 179120 119400
rect 179380 119380 179620 119400
rect 179880 119380 180120 119400
rect 180380 119380 180620 119400
rect 180880 119380 181120 119400
rect 181380 119380 182120 119400
rect 182380 119380 182620 119400
rect 182880 119380 183120 119400
rect 183380 119380 183620 119400
rect 183880 119380 184000 119400
rect 162000 119120 162100 119380
rect 162400 119120 162600 119380
rect 162900 119120 163100 119380
rect 163400 119120 163600 119380
rect 163900 119120 164100 119380
rect 164400 119120 164600 119380
rect 164900 119120 165100 119380
rect 165400 119120 165600 119380
rect 165900 119120 166100 119380
rect 166400 119120 166600 119380
rect 166900 119120 167100 119380
rect 167400 119120 167600 119380
rect 167900 119120 168100 119380
rect 168400 119120 168600 119380
rect 168900 119120 169100 119380
rect 169400 119120 169600 119380
rect 169900 119120 170100 119380
rect 170400 119120 170600 119380
rect 170900 119120 171100 119380
rect 171400 119120 171600 119380
rect 171900 119120 172100 119380
rect 172400 119120 172600 119380
rect 172900 119120 173100 119380
rect 173400 119120 173600 119380
rect 173900 119120 174100 119380
rect 174400 119120 174600 119380
rect 174900 119120 175100 119380
rect 175400 119120 175600 119380
rect 175900 119120 176100 119380
rect 176400 119120 176600 119380
rect 176900 119120 177100 119380
rect 177400 119120 177600 119380
rect 177900 119120 178100 119380
rect 178400 119120 178600 119380
rect 178900 119120 179100 119380
rect 179400 119120 179600 119380
rect 179900 119120 180100 119380
rect 180400 119120 180600 119380
rect 180900 119120 181100 119380
rect 181400 119120 182100 119380
rect 182400 119120 182600 119380
rect 182900 119120 183100 119380
rect 183400 119120 183600 119380
rect 183900 119120 184000 119380
rect 162000 119100 162120 119120
rect 162380 119100 162620 119120
rect 162880 119100 163120 119120
rect 163380 119100 163620 119120
rect 163880 119100 164120 119120
rect 164380 119100 164620 119120
rect 164880 119100 165120 119120
rect 165380 119100 165620 119120
rect 165880 119100 166120 119120
rect 166380 119100 166620 119120
rect 166880 119100 167120 119120
rect 167380 119100 167620 119120
rect 167880 119100 168120 119120
rect 168380 119100 168620 119120
rect 168880 119100 169120 119120
rect 169380 119100 169620 119120
rect 169880 119100 170120 119120
rect 170380 119100 170620 119120
rect 170880 119100 171120 119120
rect 171380 119100 171620 119120
rect 171880 119100 172120 119120
rect 172380 119100 172620 119120
rect 172880 119100 173120 119120
rect 173380 119100 173620 119120
rect 173880 119100 174120 119120
rect 174380 119100 174620 119120
rect 174880 119100 175120 119120
rect 175380 119100 175620 119120
rect 175880 119100 176120 119120
rect 176380 119100 176620 119120
rect 176880 119100 177120 119120
rect 177380 119100 177620 119120
rect 177880 119100 178120 119120
rect 178380 119100 178620 119120
rect 178880 119100 179120 119120
rect 179380 119100 179620 119120
rect 179880 119100 180120 119120
rect 180380 119100 180620 119120
rect 180880 119100 181120 119120
rect 181380 119100 182120 119120
rect 182380 119100 182620 119120
rect 182880 119100 183120 119120
rect 183380 119100 183620 119120
rect 183880 119100 184000 119120
rect 162000 118900 184000 119100
rect 162000 118880 162120 118900
rect 162380 118880 162620 118900
rect 162880 118880 163120 118900
rect 163380 118880 163620 118900
rect 163880 118880 164120 118900
rect 164380 118880 164620 118900
rect 164880 118880 165120 118900
rect 165380 118880 165620 118900
rect 165880 118880 166120 118900
rect 166380 118880 166620 118900
rect 166880 118880 167120 118900
rect 167380 118880 167620 118900
rect 167880 118880 168120 118900
rect 168380 118880 168620 118900
rect 168880 118880 169120 118900
rect 169380 118880 169620 118900
rect 169880 118880 170120 118900
rect 170380 118880 170620 118900
rect 170880 118880 171120 118900
rect 171380 118880 171620 118900
rect 171880 118880 172120 118900
rect 172380 118880 172620 118900
rect 172880 118880 173120 118900
rect 173380 118880 173620 118900
rect 173880 118880 174120 118900
rect 174380 118880 174620 118900
rect 174880 118880 175120 118900
rect 175380 118880 175620 118900
rect 175880 118880 176120 118900
rect 176380 118880 176620 118900
rect 176880 118880 177120 118900
rect 177380 118880 177620 118900
rect 177880 118880 178120 118900
rect 178380 118880 178620 118900
rect 178880 118880 179120 118900
rect 179380 118880 179620 118900
rect 179880 118880 180120 118900
rect 180380 118880 180620 118900
rect 180880 118880 181120 118900
rect 181380 118880 181620 118900
rect 181880 118880 182120 118900
rect 182380 118880 182620 118900
rect 182880 118880 183120 118900
rect 183380 118880 183620 118900
rect 183880 118880 184000 118900
rect 162000 118620 162100 118880
rect 162400 118620 162600 118880
rect 162900 118620 163100 118880
rect 163400 118620 163600 118880
rect 163900 118620 164100 118880
rect 164400 118620 164600 118880
rect 164900 118620 165100 118880
rect 165400 118620 165600 118880
rect 165900 118620 166100 118880
rect 166400 118620 166600 118880
rect 166900 118620 167100 118880
rect 167400 118620 167600 118880
rect 167900 118620 168100 118880
rect 168400 118620 168600 118880
rect 168900 118620 169100 118880
rect 169400 118620 169600 118880
rect 169900 118620 170100 118880
rect 170400 118620 170600 118880
rect 170900 118620 171100 118880
rect 171400 118620 171600 118880
rect 171900 118620 172100 118880
rect 172400 118620 172600 118880
rect 172900 118620 173100 118880
rect 173400 118620 173600 118880
rect 173900 118620 174100 118880
rect 174400 118620 174600 118880
rect 174900 118620 175100 118880
rect 175400 118620 175600 118880
rect 175900 118620 176100 118880
rect 176400 118620 176600 118880
rect 176900 118620 177100 118880
rect 177400 118620 177600 118880
rect 177900 118620 178100 118880
rect 178400 118620 178600 118880
rect 178900 118620 179100 118880
rect 179400 118620 179600 118880
rect 179900 118620 180100 118880
rect 180400 118620 180600 118880
rect 180900 118620 181100 118880
rect 181400 118620 181600 118880
rect 181900 118620 182100 118880
rect 182400 118620 182600 118880
rect 182900 118620 183100 118880
rect 183400 118620 183600 118880
rect 183900 118620 184000 118880
rect 162000 118600 162120 118620
rect 162380 118600 162620 118620
rect 162880 118600 163120 118620
rect 163380 118600 163620 118620
rect 163880 118600 164120 118620
rect 164380 118600 164620 118620
rect 164880 118600 165120 118620
rect 165380 118600 165620 118620
rect 165880 118600 166120 118620
rect 166380 118600 166620 118620
rect 166880 118600 167120 118620
rect 167380 118600 167620 118620
rect 167880 118600 168120 118620
rect 168380 118600 168620 118620
rect 168880 118600 169120 118620
rect 169380 118600 169620 118620
rect 169880 118600 170120 118620
rect 170380 118600 170620 118620
rect 170880 118600 171120 118620
rect 171380 118600 171620 118620
rect 171880 118600 172120 118620
rect 172380 118600 172620 118620
rect 172880 118600 173120 118620
rect 173380 118600 173620 118620
rect 173880 118600 174120 118620
rect 174380 118600 174620 118620
rect 174880 118600 175120 118620
rect 175380 118600 175620 118620
rect 175880 118600 176120 118620
rect 176380 118600 176620 118620
rect 176880 118600 177120 118620
rect 177380 118600 177620 118620
rect 177880 118600 178120 118620
rect 178380 118600 178620 118620
rect 178880 118600 179120 118620
rect 179380 118600 179620 118620
rect 179880 118600 180120 118620
rect 180380 118600 180620 118620
rect 180880 118600 181120 118620
rect 181380 118600 181620 118620
rect 181880 118600 182120 118620
rect 182380 118600 182620 118620
rect 182880 118600 183120 118620
rect 183380 118600 183620 118620
rect 183880 118600 184000 118620
rect 162000 118400 184000 118600
rect 162000 118380 162120 118400
rect 162380 118380 162620 118400
rect 162880 118380 163120 118400
rect 163380 118380 163620 118400
rect 163880 118380 164120 118400
rect 164380 118380 164620 118400
rect 164880 118380 165120 118400
rect 165380 118380 165620 118400
rect 165880 118380 166120 118400
rect 166380 118380 166620 118400
rect 166880 118380 167120 118400
rect 167380 118380 167620 118400
rect 167880 118380 168120 118400
rect 168380 118380 168620 118400
rect 168880 118380 169120 118400
rect 169380 118380 169620 118400
rect 169880 118380 170120 118400
rect 170380 118380 170620 118400
rect 170880 118380 171120 118400
rect 171380 118380 171620 118400
rect 171880 118380 172120 118400
rect 172380 118380 172620 118400
rect 172880 118380 173120 118400
rect 173380 118380 173620 118400
rect 173880 118380 174120 118400
rect 174380 118380 174620 118400
rect 174880 118380 175120 118400
rect 175380 118380 175620 118400
rect 175880 118380 176120 118400
rect 176380 118380 176620 118400
rect 176880 118380 177120 118400
rect 177380 118380 177620 118400
rect 177880 118380 178120 118400
rect 178380 118380 178620 118400
rect 178880 118380 179120 118400
rect 179380 118380 179620 118400
rect 179880 118380 180120 118400
rect 180380 118380 180620 118400
rect 180880 118380 181120 118400
rect 181380 118380 181620 118400
rect 181880 118380 182120 118400
rect 182380 118380 182620 118400
rect 182880 118380 183120 118400
rect 183380 118380 183620 118400
rect 183880 118380 184000 118400
rect 162000 118120 162100 118380
rect 162400 118120 162600 118380
rect 162900 118120 163100 118380
rect 163400 118120 163600 118380
rect 163900 118120 164100 118380
rect 164400 118120 164600 118380
rect 164900 118120 165100 118380
rect 165400 118120 165600 118380
rect 165900 118120 166100 118380
rect 166400 118120 166600 118380
rect 166900 118120 167100 118380
rect 167400 118120 167600 118380
rect 167900 118120 168100 118380
rect 168400 118120 168600 118380
rect 168900 118120 169100 118380
rect 169400 118120 169600 118380
rect 169900 118120 170100 118380
rect 170400 118120 170600 118380
rect 170900 118120 171100 118380
rect 171400 118120 171600 118380
rect 171900 118120 172100 118380
rect 172400 118120 172600 118380
rect 172900 118120 173100 118380
rect 173400 118120 173600 118380
rect 173900 118120 174100 118380
rect 174400 118120 174600 118380
rect 174900 118120 175100 118380
rect 175400 118120 175600 118380
rect 175900 118120 176100 118380
rect 176400 118120 176600 118380
rect 176900 118120 177100 118380
rect 177400 118120 177600 118380
rect 177900 118120 178100 118380
rect 178400 118120 178600 118380
rect 178900 118120 179100 118380
rect 179400 118120 179600 118380
rect 179900 118120 180100 118380
rect 180400 118120 180600 118380
rect 180900 118120 181100 118380
rect 181400 118120 181600 118380
rect 181900 118120 182100 118380
rect 182400 118120 182600 118380
rect 182900 118120 183100 118380
rect 183400 118120 183600 118380
rect 183900 118120 184000 118380
rect 162000 118100 162120 118120
rect 162380 118100 162620 118120
rect 162880 118100 163120 118120
rect 163380 118100 163620 118120
rect 163880 118100 164120 118120
rect 164380 118100 164620 118120
rect 164880 118100 165120 118120
rect 165380 118100 165620 118120
rect 165880 118100 166120 118120
rect 166380 118100 166620 118120
rect 166880 118100 167120 118120
rect 167380 118100 167620 118120
rect 167880 118100 168120 118120
rect 168380 118100 168620 118120
rect 168880 118100 169120 118120
rect 169380 118100 169620 118120
rect 169880 118100 170120 118120
rect 170380 118100 170620 118120
rect 170880 118100 171120 118120
rect 171380 118100 171620 118120
rect 171880 118100 172120 118120
rect 172380 118100 172620 118120
rect 172880 118100 173120 118120
rect 173380 118100 173620 118120
rect 173880 118100 174120 118120
rect 174380 118100 174620 118120
rect 174880 118100 175120 118120
rect 175380 118100 175620 118120
rect 175880 118100 176120 118120
rect 176380 118100 176620 118120
rect 176880 118100 177120 118120
rect 177380 118100 177620 118120
rect 177880 118100 178120 118120
rect 178380 118100 178620 118120
rect 178880 118100 179120 118120
rect 179380 118100 179620 118120
rect 179880 118100 180120 118120
rect 180380 118100 180620 118120
rect 180880 118100 181120 118120
rect 181380 118100 181620 118120
rect 181880 118100 182120 118120
rect 182380 118100 182620 118120
rect 182880 118100 183120 118120
rect 183380 118100 183620 118120
rect 183880 118100 184000 118120
rect 162000 117900 184000 118100
rect 162000 117880 162120 117900
rect 162380 117880 162620 117900
rect 162880 117880 163120 117900
rect 163380 117880 163620 117900
rect 163880 117880 164120 117900
rect 164380 117880 164620 117900
rect 164880 117880 165120 117900
rect 165380 117880 165620 117900
rect 165880 117880 166120 117900
rect 166380 117880 166620 117900
rect 166880 117880 167120 117900
rect 167380 117880 167620 117900
rect 167880 117880 168120 117900
rect 168380 117880 168620 117900
rect 168880 117880 169120 117900
rect 169380 117880 169620 117900
rect 169880 117880 170120 117900
rect 170380 117880 170620 117900
rect 170880 117880 171120 117900
rect 171380 117880 171620 117900
rect 171880 117880 172120 117900
rect 172380 117880 172620 117900
rect 172880 117880 173120 117900
rect 173380 117880 173620 117900
rect 173880 117880 174120 117900
rect 174380 117880 174620 117900
rect 174880 117880 175120 117900
rect 175380 117880 175620 117900
rect 175880 117880 176120 117900
rect 176380 117880 176620 117900
rect 176880 117880 177120 117900
rect 177380 117880 177620 117900
rect 177880 117880 178120 117900
rect 178380 117880 178620 117900
rect 178880 117880 179120 117900
rect 179380 117880 179620 117900
rect 179880 117880 180120 117900
rect 180380 117880 180620 117900
rect 180880 117880 181120 117900
rect 181380 117880 181620 117900
rect 181880 117880 182120 117900
rect 182380 117880 182620 117900
rect 182880 117880 183120 117900
rect 183380 117880 183620 117900
rect 183880 117880 184000 117900
rect 162000 117620 162100 117880
rect 162400 117620 162600 117880
rect 162900 117620 163100 117880
rect 163400 117620 163600 117880
rect 163900 117620 164100 117880
rect 164400 117620 164600 117880
rect 164900 117620 165100 117880
rect 165400 117620 165600 117880
rect 165900 117620 166100 117880
rect 166400 117620 166600 117880
rect 166900 117620 167100 117880
rect 167400 117620 167600 117880
rect 167900 117620 168100 117880
rect 168400 117620 168600 117880
rect 168900 117620 169100 117880
rect 169400 117620 169600 117880
rect 169900 117620 170100 117880
rect 170400 117620 170600 117880
rect 170900 117620 171100 117880
rect 171400 117620 171600 117880
rect 171900 117620 172100 117880
rect 172400 117620 172600 117880
rect 172900 117620 173100 117880
rect 173400 117620 173600 117880
rect 173900 117620 174100 117880
rect 174400 117620 174600 117880
rect 174900 117620 175100 117880
rect 175400 117620 175600 117880
rect 175900 117620 176100 117880
rect 176400 117620 176600 117880
rect 176900 117620 177100 117880
rect 177400 117620 177600 117880
rect 177900 117620 178100 117880
rect 178400 117620 178600 117880
rect 178900 117620 179100 117880
rect 179400 117620 179600 117880
rect 179900 117620 180100 117880
rect 180400 117620 180600 117880
rect 180900 117620 181100 117880
rect 181400 117620 181600 117880
rect 181900 117620 182100 117880
rect 182400 117620 182600 117880
rect 182900 117620 183100 117880
rect 183400 117620 183600 117880
rect 183900 117620 184000 117880
rect 162000 117600 162120 117620
rect 162380 117600 162620 117620
rect 162880 117600 163120 117620
rect 163380 117600 163620 117620
rect 163880 117600 164120 117620
rect 164380 117600 164620 117620
rect 164880 117600 165120 117620
rect 165380 117600 165620 117620
rect 165880 117600 166120 117620
rect 166380 117600 166620 117620
rect 166880 117600 167120 117620
rect 167380 117600 167620 117620
rect 167880 117600 168120 117620
rect 168380 117600 168620 117620
rect 168880 117600 169120 117620
rect 169380 117600 169620 117620
rect 169880 117600 170120 117620
rect 170380 117600 170620 117620
rect 170880 117600 171120 117620
rect 171380 117600 171620 117620
rect 171880 117600 172120 117620
rect 172380 117600 172620 117620
rect 172880 117600 173120 117620
rect 173380 117600 173620 117620
rect 173880 117600 174120 117620
rect 174380 117600 174620 117620
rect 174880 117600 175120 117620
rect 175380 117600 175620 117620
rect 175880 117600 176120 117620
rect 176380 117600 176620 117620
rect 176880 117600 177120 117620
rect 177380 117600 177620 117620
rect 177880 117600 178120 117620
rect 178380 117600 178620 117620
rect 178880 117600 179120 117620
rect 179380 117600 179620 117620
rect 179880 117600 180120 117620
rect 180380 117600 180620 117620
rect 180880 117600 181120 117620
rect 181380 117600 181620 117620
rect 181880 117600 182120 117620
rect 182380 117600 182620 117620
rect 182880 117600 183120 117620
rect 183380 117600 183620 117620
rect 183880 117600 184000 117620
rect 162000 117400 184000 117600
rect 162000 117380 162120 117400
rect 162380 117380 162620 117400
rect 162880 117380 163120 117400
rect 163380 117380 163620 117400
rect 163880 117380 164120 117400
rect 164380 117380 164620 117400
rect 164880 117380 165120 117400
rect 165380 117380 165620 117400
rect 165880 117380 166120 117400
rect 166380 117380 166620 117400
rect 166880 117380 167120 117400
rect 167380 117380 167620 117400
rect 167880 117380 168120 117400
rect 168380 117380 168620 117400
rect 168880 117380 169120 117400
rect 169380 117380 169620 117400
rect 169880 117380 170120 117400
rect 170380 117380 170620 117400
rect 170880 117380 171120 117400
rect 171380 117380 171620 117400
rect 171880 117380 172120 117400
rect 172380 117380 172620 117400
rect 172880 117380 173120 117400
rect 173380 117380 173620 117400
rect 173880 117380 174120 117400
rect 174380 117380 174620 117400
rect 174880 117380 175120 117400
rect 175380 117380 175620 117400
rect 175880 117380 176120 117400
rect 176380 117380 176620 117400
rect 176880 117380 177120 117400
rect 177380 117380 177620 117400
rect 177880 117380 178120 117400
rect 178380 117380 178620 117400
rect 178880 117380 179120 117400
rect 179380 117380 179620 117400
rect 179880 117380 180120 117400
rect 180380 117380 180620 117400
rect 180880 117380 181120 117400
rect 181380 117380 181620 117400
rect 181880 117380 182120 117400
rect 182380 117380 182620 117400
rect 182880 117380 183120 117400
rect 183380 117380 183620 117400
rect 183880 117380 184000 117400
rect 162000 117120 162100 117380
rect 162400 117120 162600 117380
rect 162900 117120 163100 117380
rect 163400 117120 163600 117380
rect 163900 117120 164100 117380
rect 164400 117120 164600 117380
rect 164900 117120 165100 117380
rect 165400 117120 165600 117380
rect 165900 117120 166100 117380
rect 166400 117120 166600 117380
rect 166900 117120 167100 117380
rect 167400 117120 167600 117380
rect 167900 117120 168100 117380
rect 168400 117120 168600 117380
rect 168900 117120 169100 117380
rect 169400 117120 169600 117380
rect 169900 117120 170100 117380
rect 170400 117120 170600 117380
rect 170900 117120 171100 117380
rect 171400 117120 171600 117380
rect 171900 117120 172100 117380
rect 172400 117120 172600 117380
rect 172900 117120 173100 117380
rect 173400 117120 173600 117380
rect 173900 117120 174100 117380
rect 174400 117120 174600 117380
rect 174900 117120 175100 117380
rect 175400 117120 175600 117380
rect 175900 117120 176100 117380
rect 176400 117120 176600 117380
rect 176900 117120 177100 117380
rect 177400 117120 177600 117380
rect 177900 117120 178100 117380
rect 178400 117120 178600 117380
rect 178900 117120 179100 117380
rect 179400 117120 179600 117380
rect 179900 117120 180100 117380
rect 180400 117120 180600 117380
rect 180900 117120 181100 117380
rect 181400 117120 181600 117380
rect 181900 117120 182100 117380
rect 182400 117120 182600 117380
rect 182900 117120 183100 117380
rect 183400 117120 183600 117380
rect 183900 117120 184000 117380
rect 162000 117100 162120 117120
rect 162380 117100 162620 117120
rect 162880 117100 163120 117120
rect 163380 117100 163620 117120
rect 163880 117100 164120 117120
rect 164380 117100 164620 117120
rect 164880 117100 165120 117120
rect 165380 117100 165620 117120
rect 165880 117100 166120 117120
rect 166380 117100 166620 117120
rect 166880 117100 167120 117120
rect 167380 117100 167620 117120
rect 167880 117100 168120 117120
rect 168380 117100 168620 117120
rect 168880 117100 169120 117120
rect 169380 117100 169620 117120
rect 169880 117100 170120 117120
rect 170380 117100 170620 117120
rect 170880 117100 171120 117120
rect 171380 117100 171620 117120
rect 171880 117100 172120 117120
rect 172380 117100 172620 117120
rect 172880 117100 173120 117120
rect 173380 117100 173620 117120
rect 173880 117100 174120 117120
rect 174380 117100 174620 117120
rect 174880 117100 175120 117120
rect 175380 117100 175620 117120
rect 175880 117100 176120 117120
rect 176380 117100 176620 117120
rect 176880 117100 177120 117120
rect 177380 117100 177620 117120
rect 177880 117100 178120 117120
rect 178380 117100 178620 117120
rect 178880 117100 179120 117120
rect 179380 117100 179620 117120
rect 179880 117100 180120 117120
rect 180380 117100 180620 117120
rect 180880 117100 181120 117120
rect 181380 117100 181620 117120
rect 181880 117100 182120 117120
rect 182380 117100 182620 117120
rect 182880 117100 183120 117120
rect 183380 117100 183620 117120
rect 183880 117100 184000 117120
rect 162000 116900 184000 117100
rect 162000 116880 162120 116900
rect 162380 116880 162620 116900
rect 162880 116880 163120 116900
rect 163380 116880 163620 116900
rect 163880 116880 164120 116900
rect 164380 116880 164620 116900
rect 164880 116880 165120 116900
rect 165380 116880 165620 116900
rect 165880 116880 166120 116900
rect 166380 116880 166620 116900
rect 166880 116880 167120 116900
rect 167380 116880 167620 116900
rect 167880 116880 168120 116900
rect 168380 116880 168620 116900
rect 168880 116880 169120 116900
rect 169380 116880 169620 116900
rect 169880 116880 170120 116900
rect 170380 116880 170620 116900
rect 170880 116880 171120 116900
rect 171380 116880 171620 116900
rect 171880 116880 172120 116900
rect 172380 116880 172620 116900
rect 172880 116880 173120 116900
rect 173380 116880 173620 116900
rect 173880 116880 174120 116900
rect 174380 116880 174620 116900
rect 174880 116880 175120 116900
rect 175380 116880 175620 116900
rect 175880 116880 176120 116900
rect 176380 116880 176620 116900
rect 176880 116880 177120 116900
rect 177380 116880 177620 116900
rect 177880 116880 178120 116900
rect 178380 116880 178620 116900
rect 178880 116880 179120 116900
rect 179380 116880 179620 116900
rect 179880 116880 180120 116900
rect 180380 116880 180620 116900
rect 180880 116880 181120 116900
rect 181380 116880 181620 116900
rect 181880 116880 182120 116900
rect 182380 116880 182620 116900
rect 182880 116880 183120 116900
rect 183380 116880 183620 116900
rect 183880 116880 184000 116900
rect 162000 116620 162100 116880
rect 162400 116620 162600 116880
rect 162900 116620 163100 116880
rect 163400 116620 163600 116880
rect 163900 116620 164100 116880
rect 164400 116620 164600 116880
rect 164900 116620 165100 116880
rect 165400 116620 165600 116880
rect 165900 116620 166100 116880
rect 166400 116620 166600 116880
rect 166900 116620 167100 116880
rect 167400 116620 167600 116880
rect 167900 116620 168100 116880
rect 168400 116620 168600 116880
rect 168900 116620 169100 116880
rect 169400 116620 169600 116880
rect 169900 116620 170100 116880
rect 170400 116620 170600 116880
rect 170900 116620 171100 116880
rect 171400 116620 171600 116880
rect 171900 116620 172100 116880
rect 172400 116620 172600 116880
rect 172900 116620 173100 116880
rect 173400 116620 173600 116880
rect 173900 116620 174100 116880
rect 174400 116620 174600 116880
rect 174900 116620 175100 116880
rect 175400 116620 175600 116880
rect 175900 116620 176100 116880
rect 176400 116620 176600 116880
rect 176900 116620 177100 116880
rect 177400 116620 177600 116880
rect 177900 116620 178100 116880
rect 178400 116620 178600 116880
rect 178900 116620 179100 116880
rect 179400 116620 179600 116880
rect 179900 116620 180100 116880
rect 180400 116620 180600 116880
rect 180900 116620 181100 116880
rect 181400 116620 181600 116880
rect 181900 116620 182100 116880
rect 182400 116620 182600 116880
rect 182900 116620 183100 116880
rect 183400 116620 183600 116880
rect 183900 116620 184000 116880
rect 162000 116600 162120 116620
rect 162380 116600 162620 116620
rect 162880 116600 163120 116620
rect 163380 116600 163620 116620
rect 163880 116600 164120 116620
rect 164380 116600 164620 116620
rect 164880 116600 165120 116620
rect 165380 116600 165620 116620
rect 165880 116600 166120 116620
rect 166380 116600 166620 116620
rect 166880 116600 167120 116620
rect 167380 116600 167620 116620
rect 167880 116600 168120 116620
rect 168380 116600 168620 116620
rect 168880 116600 169120 116620
rect 169380 116600 169620 116620
rect 169880 116600 170120 116620
rect 170380 116600 170620 116620
rect 170880 116600 171120 116620
rect 171380 116600 171620 116620
rect 171880 116600 172120 116620
rect 172380 116600 172620 116620
rect 172880 116600 173120 116620
rect 173380 116600 173620 116620
rect 173880 116600 174120 116620
rect 174380 116600 174620 116620
rect 174880 116600 175120 116620
rect 175380 116600 175620 116620
rect 175880 116600 176120 116620
rect 176380 116600 176620 116620
rect 176880 116600 177120 116620
rect 177380 116600 177620 116620
rect 177880 116600 178120 116620
rect 178380 116600 178620 116620
rect 178880 116600 179120 116620
rect 179380 116600 179620 116620
rect 179880 116600 180120 116620
rect 180380 116600 180620 116620
rect 180880 116600 181120 116620
rect 181380 116600 181620 116620
rect 181880 116600 182120 116620
rect 182380 116600 182620 116620
rect 182880 116600 183120 116620
rect 183380 116600 183620 116620
rect 183880 116600 184000 116620
rect 162000 116400 184000 116600
rect 162000 116380 162120 116400
rect 162380 116380 162620 116400
rect 162880 116380 163120 116400
rect 163380 116380 163620 116400
rect 163880 116380 164120 116400
rect 164380 116380 164620 116400
rect 164880 116380 165120 116400
rect 165380 116380 165620 116400
rect 165880 116380 166120 116400
rect 166380 116380 166620 116400
rect 166880 116380 167120 116400
rect 167380 116380 167620 116400
rect 167880 116380 168120 116400
rect 168380 116380 168620 116400
rect 168880 116380 169120 116400
rect 169380 116380 169620 116400
rect 169880 116380 170120 116400
rect 170380 116380 170620 116400
rect 170880 116380 171120 116400
rect 171380 116380 171620 116400
rect 171880 116380 172120 116400
rect 172380 116380 172620 116400
rect 172880 116380 173120 116400
rect 173380 116380 173620 116400
rect 173880 116380 174120 116400
rect 174380 116380 174620 116400
rect 174880 116380 175120 116400
rect 175380 116380 175620 116400
rect 175880 116380 176120 116400
rect 176380 116380 176620 116400
rect 176880 116380 177120 116400
rect 177380 116380 177620 116400
rect 177880 116380 178120 116400
rect 178380 116380 178620 116400
rect 178880 116380 179120 116400
rect 179380 116380 179620 116400
rect 179880 116380 180120 116400
rect 180380 116380 180620 116400
rect 180880 116380 181120 116400
rect 181380 116380 181620 116400
rect 181880 116380 182120 116400
rect 182380 116380 182620 116400
rect 182880 116380 183120 116400
rect 183380 116380 183620 116400
rect 183880 116380 184000 116400
rect 162000 116120 162100 116380
rect 162400 116120 162600 116380
rect 162900 116120 163100 116380
rect 163400 116120 163600 116380
rect 163900 116120 164100 116380
rect 164400 116120 164600 116380
rect 164900 116120 165100 116380
rect 165400 116120 165600 116380
rect 165900 116120 166100 116380
rect 166400 116120 166600 116380
rect 166900 116120 167100 116380
rect 167400 116120 167600 116380
rect 167900 116120 168100 116380
rect 168400 116120 168600 116380
rect 168900 116120 169100 116380
rect 169400 116120 169600 116380
rect 169900 116120 170100 116380
rect 170400 116120 170600 116380
rect 170900 116120 171100 116380
rect 171400 116120 171600 116380
rect 171900 116120 172100 116380
rect 172400 116120 172600 116380
rect 172900 116120 173100 116380
rect 173400 116120 173600 116380
rect 173900 116120 174100 116380
rect 174400 116120 174600 116380
rect 174900 116120 175100 116380
rect 175400 116120 175600 116380
rect 175900 116120 176100 116380
rect 176400 116120 176600 116380
rect 176900 116120 177100 116380
rect 177400 116120 177600 116380
rect 177900 116120 178100 116380
rect 178400 116120 178600 116380
rect 178900 116120 179100 116380
rect 179400 116120 179600 116380
rect 179900 116120 180100 116380
rect 180400 116120 180600 116380
rect 180900 116120 181100 116380
rect 181400 116120 181600 116380
rect 181900 116120 182100 116380
rect 182400 116120 182600 116380
rect 182900 116120 183100 116380
rect 183400 116120 183600 116380
rect 183900 116120 184000 116380
rect 162000 116100 162120 116120
rect 162380 116100 162620 116120
rect 162880 116100 163120 116120
rect 163380 116100 163620 116120
rect 163880 116100 164120 116120
rect 164380 116100 164620 116120
rect 164880 116100 165120 116120
rect 165380 116100 165620 116120
rect 165880 116100 166120 116120
rect 166380 116100 166620 116120
rect 166880 116100 167120 116120
rect 167380 116100 167620 116120
rect 167880 116100 168120 116120
rect 168380 116100 168620 116120
rect 168880 116100 169120 116120
rect 169380 116100 169620 116120
rect 169880 116100 170120 116120
rect 170380 116100 170620 116120
rect 170880 116100 171120 116120
rect 171380 116100 171620 116120
rect 171880 116100 172120 116120
rect 172380 116100 172620 116120
rect 172880 116100 173120 116120
rect 173380 116100 173620 116120
rect 173880 116100 174120 116120
rect 174380 116100 174620 116120
rect 174880 116100 175120 116120
rect 175380 116100 175620 116120
rect 175880 116100 176120 116120
rect 176380 116100 176620 116120
rect 176880 116100 177120 116120
rect 177380 116100 177620 116120
rect 177880 116100 178120 116120
rect 178380 116100 178620 116120
rect 178880 116100 179120 116120
rect 179380 116100 179620 116120
rect 179880 116100 180120 116120
rect 180380 116100 180620 116120
rect 180880 116100 181120 116120
rect 181380 116100 181620 116120
rect 181880 116100 182120 116120
rect 182380 116100 182620 116120
rect 182880 116100 183120 116120
rect 183380 116100 183620 116120
rect 183880 116100 184000 116120
rect 162000 115900 184000 116100
rect 162000 115880 162120 115900
rect 162380 115880 162620 115900
rect 162880 115880 163120 115900
rect 163380 115880 163620 115900
rect 163880 115880 164120 115900
rect 164380 115880 164620 115900
rect 164880 115880 165120 115900
rect 165380 115880 165620 115900
rect 165880 115880 166120 115900
rect 166380 115880 166620 115900
rect 166880 115880 167120 115900
rect 167380 115880 167620 115900
rect 167880 115880 168120 115900
rect 168380 115880 168620 115900
rect 168880 115880 169120 115900
rect 169380 115880 169620 115900
rect 169880 115880 170120 115900
rect 170380 115880 170620 115900
rect 170880 115880 171120 115900
rect 171380 115880 171620 115900
rect 171880 115880 172120 115900
rect 172380 115880 172620 115900
rect 172880 115880 173120 115900
rect 173380 115880 173620 115900
rect 173880 115880 174120 115900
rect 174380 115880 174620 115900
rect 174880 115880 175120 115900
rect 175380 115880 175620 115900
rect 175880 115880 176120 115900
rect 176380 115880 176620 115900
rect 176880 115880 177120 115900
rect 177380 115880 177620 115900
rect 177880 115880 178120 115900
rect 178380 115880 178620 115900
rect 178880 115880 179120 115900
rect 179380 115880 179620 115900
rect 179880 115880 180120 115900
rect 180380 115880 180620 115900
rect 180880 115880 181120 115900
rect 181380 115880 181620 115900
rect 181880 115880 182120 115900
rect 182380 115880 182620 115900
rect 182880 115880 183120 115900
rect 183380 115880 183620 115900
rect 183880 115880 184000 115900
rect 162000 115620 162100 115880
rect 162400 115620 162600 115880
rect 162900 115620 163100 115880
rect 163400 115620 163600 115880
rect 163900 115620 164100 115880
rect 164400 115620 164600 115880
rect 164900 115620 165100 115880
rect 165400 115620 165600 115880
rect 165900 115620 166100 115880
rect 166400 115620 166600 115880
rect 166900 115620 167100 115880
rect 167400 115620 167600 115880
rect 167900 115620 168100 115880
rect 168400 115620 168600 115880
rect 168900 115620 169100 115880
rect 169400 115620 169600 115880
rect 169900 115620 170100 115880
rect 170400 115620 170600 115880
rect 170900 115620 171100 115880
rect 171400 115620 171600 115880
rect 171900 115620 172100 115880
rect 172400 115620 172600 115880
rect 172900 115620 173100 115880
rect 173400 115620 173600 115880
rect 173900 115620 174100 115880
rect 174400 115620 174600 115880
rect 174900 115620 175100 115880
rect 175400 115620 175600 115880
rect 175900 115620 176100 115880
rect 176400 115620 176600 115880
rect 176900 115620 177100 115880
rect 177400 115620 177600 115880
rect 177900 115620 178100 115880
rect 178400 115620 178600 115880
rect 178900 115620 179100 115880
rect 179400 115620 179600 115880
rect 179900 115620 180100 115880
rect 180400 115620 180600 115880
rect 180900 115620 181100 115880
rect 181400 115620 181600 115880
rect 181900 115620 182100 115880
rect 182400 115620 182600 115880
rect 182900 115620 183100 115880
rect 183400 115620 183600 115880
rect 183900 115620 184000 115880
rect 162000 115600 162120 115620
rect 162380 115600 162620 115620
rect 162880 115600 163120 115620
rect 163380 115600 163620 115620
rect 163880 115600 164120 115620
rect 164380 115600 164620 115620
rect 164880 115600 165120 115620
rect 165380 115600 165620 115620
rect 165880 115600 166120 115620
rect 166380 115600 166620 115620
rect 166880 115600 167120 115620
rect 167380 115600 167620 115620
rect 167880 115600 168120 115620
rect 168380 115600 168620 115620
rect 168880 115600 169120 115620
rect 169380 115600 169620 115620
rect 169880 115600 170120 115620
rect 170380 115600 170620 115620
rect 170880 115600 171120 115620
rect 171380 115600 171620 115620
rect 171880 115600 172120 115620
rect 172380 115600 172620 115620
rect 172880 115600 173120 115620
rect 173380 115600 173620 115620
rect 173880 115600 174120 115620
rect 174380 115600 174620 115620
rect 174880 115600 175120 115620
rect 175380 115600 175620 115620
rect 175880 115600 176120 115620
rect 176380 115600 176620 115620
rect 176880 115600 177120 115620
rect 177380 115600 177620 115620
rect 177880 115600 178120 115620
rect 178380 115600 178620 115620
rect 178880 115600 179120 115620
rect 179380 115600 179620 115620
rect 179880 115600 180120 115620
rect 180380 115600 180620 115620
rect 180880 115600 181120 115620
rect 181380 115600 181620 115620
rect 181880 115600 182120 115620
rect 182380 115600 182620 115620
rect 182880 115600 183120 115620
rect 183380 115600 183620 115620
rect 183880 115600 184000 115620
rect 162000 115400 184000 115600
rect 162000 115380 162120 115400
rect 162380 115380 162620 115400
rect 162880 115380 163120 115400
rect 163380 115380 163620 115400
rect 163880 115380 164120 115400
rect 164380 115380 164620 115400
rect 164880 115380 165120 115400
rect 165380 115380 165620 115400
rect 165880 115380 166120 115400
rect 166380 115380 166620 115400
rect 166880 115380 167120 115400
rect 167380 115380 167620 115400
rect 167880 115380 168120 115400
rect 168380 115380 168620 115400
rect 168880 115380 169120 115400
rect 169380 115380 169620 115400
rect 169880 115380 170120 115400
rect 170380 115380 170620 115400
rect 170880 115380 171120 115400
rect 171380 115380 171620 115400
rect 171880 115380 172120 115400
rect 172380 115380 172620 115400
rect 172880 115380 173120 115400
rect 173380 115380 173620 115400
rect 173880 115380 174120 115400
rect 174380 115380 174620 115400
rect 174880 115380 175120 115400
rect 175380 115380 175620 115400
rect 175880 115380 176120 115400
rect 176380 115380 176620 115400
rect 176880 115380 177120 115400
rect 177380 115380 177620 115400
rect 177880 115380 178120 115400
rect 178380 115380 178620 115400
rect 178880 115380 179120 115400
rect 179380 115380 179620 115400
rect 179880 115380 180120 115400
rect 180380 115380 180620 115400
rect 180880 115380 181120 115400
rect 181380 115380 181620 115400
rect 181880 115380 182120 115400
rect 182380 115380 182620 115400
rect 182880 115380 183120 115400
rect 183380 115380 183620 115400
rect 183880 115380 184000 115400
rect 162000 115120 162100 115380
rect 162400 115120 162600 115380
rect 162900 115120 163100 115380
rect 163400 115120 163600 115380
rect 163900 115120 164100 115380
rect 164400 115120 164600 115380
rect 164900 115120 165100 115380
rect 165400 115120 165600 115380
rect 165900 115120 166100 115380
rect 166400 115120 166600 115380
rect 166900 115120 167100 115380
rect 167400 115120 167600 115380
rect 167900 115120 168100 115380
rect 168400 115120 168600 115380
rect 168900 115120 169100 115380
rect 169400 115120 169600 115380
rect 169900 115120 170100 115380
rect 170400 115120 170600 115380
rect 170900 115120 171100 115380
rect 171400 115120 171600 115380
rect 171900 115120 172100 115380
rect 172400 115120 172600 115380
rect 172900 115120 173100 115380
rect 173400 115120 173600 115380
rect 173900 115120 174100 115380
rect 174400 115120 174600 115380
rect 174900 115120 175100 115380
rect 175400 115120 175600 115380
rect 175900 115120 176100 115380
rect 176400 115120 176600 115380
rect 176900 115120 177100 115380
rect 177400 115120 177600 115380
rect 177900 115120 178100 115380
rect 178400 115120 178600 115380
rect 178900 115120 179100 115380
rect 179400 115120 179600 115380
rect 179900 115120 180100 115380
rect 180400 115120 180600 115380
rect 180900 115120 181100 115380
rect 181400 115120 181600 115380
rect 181900 115120 182100 115380
rect 182400 115120 182600 115380
rect 182900 115120 183100 115380
rect 183400 115120 183600 115380
rect 183900 115120 184000 115380
rect 162000 115100 162120 115120
rect 162380 115100 162620 115120
rect 162880 115100 163120 115120
rect 163380 115100 163620 115120
rect 163880 115100 164120 115120
rect 164380 115100 164620 115120
rect 164880 115100 165120 115120
rect 165380 115100 165620 115120
rect 165880 115100 166120 115120
rect 166380 115100 166620 115120
rect 166880 115100 167120 115120
rect 167380 115100 167620 115120
rect 167880 115100 168120 115120
rect 168380 115100 168620 115120
rect 168880 115100 169120 115120
rect 169380 115100 169620 115120
rect 169880 115100 170120 115120
rect 170380 115100 170620 115120
rect 170880 115100 171120 115120
rect 171380 115100 171620 115120
rect 171880 115100 172120 115120
rect 172380 115100 172620 115120
rect 172880 115100 173120 115120
rect 173380 115100 173620 115120
rect 173880 115100 174120 115120
rect 174380 115100 174620 115120
rect 174880 115100 175120 115120
rect 175380 115100 175620 115120
rect 175880 115100 176120 115120
rect 176380 115100 176620 115120
rect 176880 115100 177120 115120
rect 177380 115100 177620 115120
rect 177880 115100 178120 115120
rect 178380 115100 178620 115120
rect 178880 115100 179120 115120
rect 179380 115100 179620 115120
rect 179880 115100 180120 115120
rect 180380 115100 180620 115120
rect 180880 115100 181120 115120
rect 181380 115100 181620 115120
rect 181880 115100 182120 115120
rect 182380 115100 182620 115120
rect 182880 115100 183120 115120
rect 183380 115100 183620 115120
rect 183880 115100 184000 115120
rect 162000 114900 184000 115100
rect 162000 114880 162120 114900
rect 162380 114880 162620 114900
rect 162880 114880 163120 114900
rect 163380 114880 163620 114900
rect 163880 114880 164120 114900
rect 164380 114880 164620 114900
rect 164880 114880 165120 114900
rect 165380 114880 165620 114900
rect 165880 114880 166120 114900
rect 166380 114880 166620 114900
rect 166880 114880 167120 114900
rect 167380 114880 167620 114900
rect 167880 114880 168120 114900
rect 168380 114880 168620 114900
rect 168880 114880 169120 114900
rect 169380 114880 169620 114900
rect 169880 114880 170120 114900
rect 170380 114880 170620 114900
rect 170880 114880 171120 114900
rect 171380 114880 171620 114900
rect 171880 114880 172120 114900
rect 172380 114880 172620 114900
rect 172880 114880 173120 114900
rect 173380 114880 173620 114900
rect 173880 114880 174120 114900
rect 174380 114880 174620 114900
rect 174880 114880 175120 114900
rect 175380 114880 175620 114900
rect 175880 114880 176120 114900
rect 176380 114880 176620 114900
rect 176880 114880 177120 114900
rect 177380 114880 177620 114900
rect 177880 114880 178120 114900
rect 178380 114880 178620 114900
rect 178880 114880 179120 114900
rect 179380 114880 179620 114900
rect 179880 114880 180120 114900
rect 180380 114880 180620 114900
rect 180880 114880 181120 114900
rect 181380 114880 181620 114900
rect 181880 114880 182120 114900
rect 182380 114880 182620 114900
rect 182880 114880 183120 114900
rect 183380 114880 183620 114900
rect 183880 114880 184000 114900
rect 162000 114620 162100 114880
rect 162400 114620 162600 114880
rect 162900 114620 163100 114880
rect 163400 114620 163600 114880
rect 163900 114620 164100 114880
rect 164400 114620 164600 114880
rect 164900 114620 165100 114880
rect 165400 114620 165600 114880
rect 165900 114620 166100 114880
rect 166400 114620 166600 114880
rect 166900 114620 167100 114880
rect 167400 114620 167600 114880
rect 167900 114620 168100 114880
rect 168400 114620 168600 114880
rect 168900 114620 169100 114880
rect 169400 114620 169600 114880
rect 169900 114620 170100 114880
rect 170400 114620 170600 114880
rect 170900 114620 171100 114880
rect 171400 114620 171600 114880
rect 171900 114620 172100 114880
rect 172400 114620 172600 114880
rect 172900 114620 173100 114880
rect 173400 114620 173600 114880
rect 173900 114620 174100 114880
rect 174400 114620 174600 114880
rect 174900 114620 175100 114880
rect 175400 114620 175600 114880
rect 175900 114620 176100 114880
rect 176400 114620 176600 114880
rect 176900 114620 177100 114880
rect 177400 114620 177600 114880
rect 177900 114620 178100 114880
rect 178400 114620 178600 114880
rect 178900 114620 179100 114880
rect 179400 114620 179600 114880
rect 179900 114620 180100 114880
rect 180400 114620 180600 114880
rect 180900 114620 181100 114880
rect 181400 114620 181600 114880
rect 181900 114620 182100 114880
rect 182400 114620 182600 114880
rect 182900 114620 183100 114880
rect 183400 114620 183600 114880
rect 183900 114620 184000 114880
rect 162000 114600 162120 114620
rect 162380 114600 162620 114620
rect 162880 114600 163120 114620
rect 163380 114600 163620 114620
rect 163880 114600 164120 114620
rect 164380 114600 164620 114620
rect 164880 114600 165120 114620
rect 165380 114600 165620 114620
rect 165880 114600 166120 114620
rect 166380 114600 166620 114620
rect 166880 114600 167120 114620
rect 167380 114600 167620 114620
rect 167880 114600 168120 114620
rect 168380 114600 168620 114620
rect 168880 114600 169120 114620
rect 169380 114600 169620 114620
rect 169880 114600 170120 114620
rect 170380 114600 170620 114620
rect 170880 114600 171120 114620
rect 171380 114600 171620 114620
rect 171880 114600 172120 114620
rect 172380 114600 172620 114620
rect 172880 114600 173120 114620
rect 173380 114600 173620 114620
rect 173880 114600 174120 114620
rect 174380 114600 174620 114620
rect 174880 114600 175120 114620
rect 175380 114600 175620 114620
rect 175880 114600 176120 114620
rect 176380 114600 176620 114620
rect 176880 114600 177120 114620
rect 177380 114600 177620 114620
rect 177880 114600 178120 114620
rect 178380 114600 178620 114620
rect 178880 114600 179120 114620
rect 179380 114600 179620 114620
rect 179880 114600 180120 114620
rect 180380 114600 180620 114620
rect 180880 114600 181120 114620
rect 181380 114600 181620 114620
rect 181880 114600 182120 114620
rect 182380 114600 182620 114620
rect 182880 114600 183120 114620
rect 183380 114600 183620 114620
rect 183880 114600 184000 114620
rect 162000 114400 184000 114600
rect 162000 114380 162120 114400
rect 162380 114380 162620 114400
rect 162880 114380 163120 114400
rect 163380 114380 163620 114400
rect 163880 114380 164120 114400
rect 164380 114380 164620 114400
rect 164880 114380 165120 114400
rect 165380 114380 165620 114400
rect 165880 114380 166120 114400
rect 166380 114380 166620 114400
rect 166880 114380 167120 114400
rect 167380 114380 167620 114400
rect 167880 114380 168120 114400
rect 168380 114380 168620 114400
rect 168880 114380 169120 114400
rect 169380 114380 169620 114400
rect 169880 114380 170120 114400
rect 170380 114380 170620 114400
rect 170880 114380 171120 114400
rect 171380 114380 171620 114400
rect 171880 114380 172120 114400
rect 172380 114380 172620 114400
rect 172880 114380 173120 114400
rect 173380 114380 173620 114400
rect 173880 114380 174120 114400
rect 174380 114380 174620 114400
rect 174880 114380 175120 114400
rect 175380 114380 175620 114400
rect 175880 114380 176120 114400
rect 176380 114380 176620 114400
rect 176880 114380 177120 114400
rect 177380 114380 177620 114400
rect 177880 114380 178120 114400
rect 178380 114380 178620 114400
rect 178880 114380 179120 114400
rect 179380 114380 179620 114400
rect 179880 114380 180120 114400
rect 180380 114380 180620 114400
rect 180880 114380 181120 114400
rect 181380 114380 181620 114400
rect 181880 114380 182120 114400
rect 182380 114380 182620 114400
rect 182880 114380 183120 114400
rect 183380 114380 183620 114400
rect 183880 114380 184000 114400
rect 162000 114120 162100 114380
rect 162400 114120 162600 114380
rect 162900 114120 163100 114380
rect 163400 114120 163600 114380
rect 163900 114120 164100 114380
rect 164400 114120 164600 114380
rect 164900 114120 165100 114380
rect 165400 114120 165600 114380
rect 165900 114120 166100 114380
rect 166400 114120 166600 114380
rect 166900 114120 167100 114380
rect 167400 114120 167600 114380
rect 167900 114120 168100 114380
rect 168400 114120 168600 114380
rect 168900 114120 169100 114380
rect 169400 114120 169600 114380
rect 169900 114120 170100 114380
rect 170400 114120 170600 114380
rect 170900 114120 171100 114380
rect 171400 114120 171600 114380
rect 171900 114120 172100 114380
rect 172400 114120 172600 114380
rect 172900 114120 173100 114380
rect 173400 114120 173600 114380
rect 173900 114120 174100 114380
rect 174400 114120 174600 114380
rect 174900 114120 175100 114380
rect 175400 114120 175600 114380
rect 175900 114120 176100 114380
rect 176400 114120 176600 114380
rect 176900 114120 177100 114380
rect 177400 114120 177600 114380
rect 177900 114120 178100 114380
rect 178400 114120 178600 114380
rect 178900 114120 179100 114380
rect 179400 114120 179600 114380
rect 179900 114120 180100 114380
rect 180400 114120 180600 114380
rect 180900 114120 181100 114380
rect 181400 114120 181600 114380
rect 181900 114120 182100 114380
rect 182400 114120 182600 114380
rect 182900 114120 183100 114380
rect 183400 114120 183600 114380
rect 183900 114120 184000 114380
rect 162000 114100 162120 114120
rect 162380 114100 162620 114120
rect 162880 114100 163120 114120
rect 163380 114100 163620 114120
rect 163880 114100 164120 114120
rect 164380 114100 164620 114120
rect 164880 114100 165120 114120
rect 165380 114100 165620 114120
rect 165880 114100 166120 114120
rect 166380 114100 166620 114120
rect 166880 114100 167120 114120
rect 167380 114100 167620 114120
rect 167880 114100 168120 114120
rect 168380 114100 168620 114120
rect 168880 114100 169120 114120
rect 169380 114100 169620 114120
rect 169880 114100 170120 114120
rect 170380 114100 170620 114120
rect 170880 114100 171120 114120
rect 171380 114100 171620 114120
rect 171880 114100 172120 114120
rect 172380 114100 172620 114120
rect 172880 114100 173120 114120
rect 173380 114100 173620 114120
rect 173880 114100 174120 114120
rect 174380 114100 174620 114120
rect 174880 114100 175120 114120
rect 175380 114100 175620 114120
rect 175880 114100 176120 114120
rect 176380 114100 176620 114120
rect 176880 114100 177120 114120
rect 177380 114100 177620 114120
rect 177880 114100 178120 114120
rect 178380 114100 178620 114120
rect 178880 114100 179120 114120
rect 179380 114100 179620 114120
rect 179880 114100 180120 114120
rect 180380 114100 180620 114120
rect 180880 114100 181120 114120
rect 181380 114100 181620 114120
rect 181880 114100 182120 114120
rect 182380 114100 182620 114120
rect 182880 114100 183120 114120
rect 183380 114100 183620 114120
rect 183880 114100 184000 114120
rect 162000 114000 184000 114100
rect 214000 121900 234000 122000
rect 214000 121880 214120 121900
rect 214380 121880 214620 121900
rect 214880 121880 215120 121900
rect 215380 121880 215620 121900
rect 215880 121880 216120 121900
rect 216380 121880 216620 121900
rect 216880 121880 217120 121900
rect 217380 121880 217620 121900
rect 217880 121880 218120 121900
rect 218380 121880 218620 121900
rect 218880 121880 219120 121900
rect 219380 121880 219620 121900
rect 219880 121880 220120 121900
rect 220380 121880 220620 121900
rect 220880 121880 221120 121900
rect 221380 121880 221620 121900
rect 221880 121880 222120 121900
rect 222380 121880 222700 121900
rect 214000 121620 214100 121880
rect 214400 121620 214600 121880
rect 214900 121620 215100 121880
rect 215400 121620 215600 121880
rect 215900 121620 216100 121880
rect 216400 121620 216600 121880
rect 216900 121620 217100 121880
rect 217400 121620 217600 121880
rect 217900 121620 218100 121880
rect 218400 121620 218600 121880
rect 218900 121620 219100 121880
rect 219400 121620 219600 121880
rect 219900 121620 220100 121880
rect 220400 121620 220600 121880
rect 220900 121620 221100 121880
rect 221400 121620 221600 121880
rect 221900 121620 222100 121880
rect 222400 121620 222700 121880
rect 214000 121600 214120 121620
rect 214380 121600 214620 121620
rect 214880 121600 215120 121620
rect 215380 121600 215620 121620
rect 215880 121600 216120 121620
rect 216380 121600 216620 121620
rect 216880 121600 217120 121620
rect 217380 121600 217620 121620
rect 217880 121600 218120 121620
rect 218380 121600 218620 121620
rect 218880 121600 219120 121620
rect 219380 121600 219620 121620
rect 219880 121600 220120 121620
rect 220380 121600 220620 121620
rect 220880 121600 221120 121620
rect 221380 121600 221620 121620
rect 221880 121600 222120 121620
rect 222380 121600 222700 121620
rect 214000 121400 222700 121600
rect 214000 121380 214120 121400
rect 214380 121380 214620 121400
rect 214880 121380 215120 121400
rect 215380 121380 215620 121400
rect 215880 121380 216120 121400
rect 216380 121380 216620 121400
rect 216880 121380 217120 121400
rect 217380 121380 217620 121400
rect 217880 121380 218120 121400
rect 218380 121380 218620 121400
rect 218880 121380 219120 121400
rect 219380 121380 219620 121400
rect 219880 121380 220120 121400
rect 220380 121380 220620 121400
rect 220880 121380 221120 121400
rect 221380 121380 221620 121400
rect 221880 121380 222120 121400
rect 222380 121380 222700 121400
rect 214000 121120 214100 121380
rect 214400 121120 214600 121380
rect 214900 121120 215100 121380
rect 215400 121120 215600 121380
rect 215900 121120 216100 121380
rect 216400 121120 216600 121380
rect 216900 121120 217100 121380
rect 217400 121120 217600 121380
rect 217900 121120 218100 121380
rect 218400 121120 218600 121380
rect 218900 121120 219100 121380
rect 219400 121120 219600 121380
rect 219900 121120 220100 121380
rect 220400 121120 220600 121380
rect 220900 121120 221100 121380
rect 221400 121120 221600 121380
rect 221900 121120 222100 121380
rect 222400 121120 222700 121380
rect 214000 121100 214120 121120
rect 214380 121100 214620 121120
rect 214880 121100 215120 121120
rect 215380 121100 215620 121120
rect 215880 121100 216120 121120
rect 216380 121100 216620 121120
rect 216880 121100 217120 121120
rect 217380 121100 217620 121120
rect 217880 121100 218120 121120
rect 218380 121100 218620 121120
rect 218880 121100 219120 121120
rect 219380 121100 219620 121120
rect 219880 121100 220120 121120
rect 220380 121100 220620 121120
rect 220880 121100 221120 121120
rect 221380 121100 221620 121120
rect 221880 121100 222120 121120
rect 222380 121100 222700 121120
rect 214000 120900 222700 121100
rect 214000 120880 214120 120900
rect 214380 120880 214620 120900
rect 214880 120880 215120 120900
rect 215380 120880 215620 120900
rect 215880 120880 216120 120900
rect 216380 120880 216620 120900
rect 216880 120880 217120 120900
rect 217380 120880 217620 120900
rect 217880 120880 218120 120900
rect 218380 120880 218620 120900
rect 218880 120880 219120 120900
rect 219380 120880 219620 120900
rect 219880 120880 220120 120900
rect 220380 120880 220620 120900
rect 220880 120880 221120 120900
rect 221380 120880 221620 120900
rect 221880 120880 222120 120900
rect 222380 120880 222700 120900
rect 214000 120620 214100 120880
rect 214400 120620 214600 120880
rect 214900 120620 215100 120880
rect 215400 120620 215600 120880
rect 215900 120620 216100 120880
rect 216400 120620 216600 120880
rect 216900 120620 217100 120880
rect 217400 120620 217600 120880
rect 217900 120620 218100 120880
rect 218400 120620 218600 120880
rect 218900 120620 219100 120880
rect 219400 120620 219600 120880
rect 219900 120620 220100 120880
rect 220400 120620 220600 120880
rect 220900 120620 221100 120880
rect 221400 120620 221600 120880
rect 221900 120620 222100 120880
rect 222400 120620 222700 120880
rect 214000 120600 214120 120620
rect 214380 120600 214620 120620
rect 214880 120600 215120 120620
rect 215380 120600 215620 120620
rect 215880 120600 216120 120620
rect 216380 120600 216620 120620
rect 216880 120600 217120 120620
rect 217380 120600 217620 120620
rect 217880 120600 218120 120620
rect 218380 120600 218620 120620
rect 218880 120600 219120 120620
rect 219380 120600 219620 120620
rect 219880 120600 220120 120620
rect 220380 120600 220620 120620
rect 220880 120600 221120 120620
rect 221380 120600 221620 120620
rect 221880 120600 222120 120620
rect 222380 120600 222700 120620
rect 214000 120400 222700 120600
rect 214000 120380 214120 120400
rect 214380 120380 214620 120400
rect 214880 120380 215120 120400
rect 215380 120380 215620 120400
rect 215880 120380 216120 120400
rect 216380 120380 216620 120400
rect 216880 120380 217120 120400
rect 217380 120380 217620 120400
rect 217880 120380 218120 120400
rect 218380 120380 218620 120400
rect 218880 120380 219120 120400
rect 219380 120380 219620 120400
rect 219880 120380 220120 120400
rect 220380 120380 220620 120400
rect 220880 120380 221120 120400
rect 221380 120380 221620 120400
rect 221880 120380 222120 120400
rect 222380 120380 222700 120400
rect 214000 120120 214100 120380
rect 214400 120120 214600 120380
rect 214900 120120 215100 120380
rect 215400 120120 215600 120380
rect 215900 120120 216100 120380
rect 216400 120120 216600 120380
rect 216900 120120 217100 120380
rect 217400 120120 217600 120380
rect 217900 120120 218100 120380
rect 218400 120120 218600 120380
rect 218900 120120 219100 120380
rect 219400 120120 219600 120380
rect 219900 120120 220100 120380
rect 220400 120120 220600 120380
rect 220900 120120 221100 120380
rect 221400 120120 221600 120380
rect 221900 120120 222100 120380
rect 222400 120120 222700 120380
rect 214000 120100 214120 120120
rect 214380 120100 214620 120120
rect 214880 120100 215120 120120
rect 215380 120100 215620 120120
rect 215880 120100 216120 120120
rect 216380 120100 216620 120120
rect 216880 120100 217120 120120
rect 217380 120100 217620 120120
rect 217880 120100 218120 120120
rect 218380 120100 218620 120120
rect 218880 120100 219120 120120
rect 219380 120100 219620 120120
rect 219880 120100 220120 120120
rect 220380 120100 220620 120120
rect 220880 120100 221120 120120
rect 221380 120100 221620 120120
rect 221880 120100 222120 120120
rect 222380 120100 222700 120120
rect 214000 119900 222700 120100
rect 214000 119880 214120 119900
rect 214380 119880 214620 119900
rect 214880 119880 215120 119900
rect 215380 119880 215620 119900
rect 215880 119880 216120 119900
rect 216380 119880 216620 119900
rect 216880 119880 217120 119900
rect 217380 119880 217620 119900
rect 217880 119880 218120 119900
rect 218380 119880 218620 119900
rect 218880 119880 219120 119900
rect 219380 119880 219620 119900
rect 219880 119880 220120 119900
rect 220380 119880 220620 119900
rect 220880 119880 221120 119900
rect 221380 119880 221620 119900
rect 221880 119880 222120 119900
rect 222380 119880 222700 119900
rect 214000 119620 214100 119880
rect 214400 119620 214600 119880
rect 214900 119620 215100 119880
rect 215400 119620 215600 119880
rect 215900 119620 216100 119880
rect 216400 119620 216600 119880
rect 216900 119620 217100 119880
rect 217400 119620 217600 119880
rect 217900 119620 218100 119880
rect 218400 119620 218600 119880
rect 218900 119620 219100 119880
rect 219400 119620 219600 119880
rect 219900 119620 220100 119880
rect 220400 119620 220600 119880
rect 220900 119620 221100 119880
rect 221400 119620 221600 119880
rect 221900 119620 222100 119880
rect 222400 119620 222700 119880
rect 214000 119600 214120 119620
rect 214380 119600 214620 119620
rect 214880 119600 215120 119620
rect 215380 119600 215620 119620
rect 215880 119600 216120 119620
rect 216380 119600 216620 119620
rect 216880 119600 217120 119620
rect 217380 119600 217620 119620
rect 217880 119600 218120 119620
rect 218380 119600 218620 119620
rect 218880 119600 219120 119620
rect 219380 119600 219620 119620
rect 219880 119600 220120 119620
rect 220380 119600 220620 119620
rect 220880 119600 221120 119620
rect 221380 119600 221620 119620
rect 221880 119600 222120 119620
rect 222380 119600 222700 119620
rect 214000 119500 222700 119600
rect 231900 121880 232120 121900
rect 232380 121880 232620 121900
rect 232880 121880 233120 121900
rect 233380 121880 233620 121900
rect 233880 121880 234000 121900
rect 231900 121620 232100 121880
rect 232400 121620 232600 121880
rect 232900 121620 233100 121880
rect 233400 121620 233600 121880
rect 233900 121620 234000 121880
rect 231900 121600 232120 121620
rect 232380 121600 232620 121620
rect 232880 121600 233120 121620
rect 233380 121600 233620 121620
rect 233880 121600 234000 121620
rect 231900 121400 234000 121600
rect 231900 121380 232120 121400
rect 232380 121380 232620 121400
rect 232880 121380 233120 121400
rect 233380 121380 233620 121400
rect 233880 121380 234000 121400
rect 231900 121120 232100 121380
rect 232400 121120 232600 121380
rect 232900 121120 233100 121380
rect 233400 121120 233600 121380
rect 233900 121120 234000 121380
rect 231900 121100 232120 121120
rect 232380 121100 232620 121120
rect 232880 121100 233120 121120
rect 233380 121100 233620 121120
rect 233880 121100 234000 121120
rect 231900 120900 234000 121100
rect 231900 120880 232120 120900
rect 232380 120880 232620 120900
rect 232880 120880 233120 120900
rect 233380 120880 233620 120900
rect 233880 120880 234000 120900
rect 231900 120620 232100 120880
rect 232400 120620 232600 120880
rect 232900 120620 233100 120880
rect 233400 120620 233600 120880
rect 233900 120620 234000 120880
rect 231900 120600 232120 120620
rect 232380 120600 232620 120620
rect 232880 120600 233120 120620
rect 233380 120600 233620 120620
rect 233880 120600 234000 120620
rect 231900 120400 234000 120600
rect 231900 120380 232120 120400
rect 232380 120380 232620 120400
rect 232880 120380 233120 120400
rect 233380 120380 233620 120400
rect 233880 120380 234000 120400
rect 231900 120120 232100 120380
rect 232400 120120 232600 120380
rect 232900 120120 233100 120380
rect 233400 120120 233600 120380
rect 233900 120120 234000 120380
rect 231900 120100 232120 120120
rect 232380 120100 232620 120120
rect 232880 120100 233120 120120
rect 233380 120100 233620 120120
rect 233880 120100 234000 120120
rect 231900 120000 234000 120100
rect 231900 119500 232000 120000
rect 214000 119400 232000 119500
rect 214000 119380 214120 119400
rect 214380 119380 214620 119400
rect 214880 119380 215120 119400
rect 215380 119380 215620 119400
rect 215880 119380 216120 119400
rect 216380 119380 216620 119400
rect 216880 119380 217120 119400
rect 217380 119380 217620 119400
rect 217880 119380 218120 119400
rect 218380 119380 218620 119400
rect 218880 119380 219120 119400
rect 219380 119380 219620 119400
rect 219880 119380 220120 119400
rect 220380 119380 220620 119400
rect 220880 119380 221120 119400
rect 221380 119380 221620 119400
rect 221880 119380 222120 119400
rect 222380 119380 222620 119400
rect 222880 119380 223120 119400
rect 223380 119380 223620 119400
rect 223880 119380 224120 119400
rect 224380 119380 224620 119400
rect 224880 119380 225120 119400
rect 225380 119380 225620 119400
rect 225880 119380 226120 119400
rect 226380 119380 226620 119400
rect 226880 119380 227120 119400
rect 227380 119380 227620 119400
rect 227880 119380 228120 119400
rect 228380 119380 228620 119400
rect 228880 119380 229120 119400
rect 229380 119380 229620 119400
rect 229880 119380 230120 119400
rect 230380 119380 230620 119400
rect 230880 119380 231120 119400
rect 231380 119380 232000 119400
rect 214000 119120 214100 119380
rect 214400 119120 214600 119380
rect 214900 119120 215100 119380
rect 215400 119120 215600 119380
rect 215900 119120 216100 119380
rect 216400 119120 216600 119380
rect 216900 119120 217100 119380
rect 217400 119120 217600 119380
rect 217900 119120 218100 119380
rect 218400 119120 218600 119380
rect 218900 119120 219100 119380
rect 219400 119120 219600 119380
rect 219900 119120 220100 119380
rect 220400 119120 220600 119380
rect 220900 119120 221100 119380
rect 221400 119120 221600 119380
rect 221900 119120 222100 119380
rect 222400 119120 222600 119380
rect 222900 119120 223100 119380
rect 223400 119120 223600 119380
rect 223900 119120 224100 119380
rect 224400 119120 224600 119380
rect 224900 119120 225100 119380
rect 225400 119120 225600 119380
rect 225900 119120 226100 119380
rect 226400 119120 226600 119380
rect 226900 119120 227100 119380
rect 227400 119120 227600 119380
rect 227900 119120 228100 119380
rect 228400 119120 228600 119380
rect 228900 119120 229100 119380
rect 229400 119120 229600 119380
rect 229900 119120 230100 119380
rect 230400 119120 230600 119380
rect 230900 119120 231100 119380
rect 231400 119120 232000 119380
rect 214000 119100 214120 119120
rect 214380 119100 214620 119120
rect 214880 119100 215120 119120
rect 215380 119100 215620 119120
rect 215880 119100 216120 119120
rect 216380 119100 216620 119120
rect 216880 119100 217120 119120
rect 217380 119100 217620 119120
rect 217880 119100 218120 119120
rect 218380 119100 218620 119120
rect 218880 119100 219120 119120
rect 219380 119100 219620 119120
rect 219880 119100 220120 119120
rect 220380 119100 220620 119120
rect 220880 119100 221120 119120
rect 221380 119100 221620 119120
rect 221880 119100 222120 119120
rect 222380 119100 222620 119120
rect 222880 119100 223120 119120
rect 223380 119100 223620 119120
rect 223880 119100 224120 119120
rect 224380 119100 224620 119120
rect 224880 119100 225120 119120
rect 225380 119100 225620 119120
rect 225880 119100 226120 119120
rect 226380 119100 226620 119120
rect 226880 119100 227120 119120
rect 227380 119100 227620 119120
rect 227880 119100 228120 119120
rect 228380 119100 228620 119120
rect 228880 119100 229120 119120
rect 229380 119100 229620 119120
rect 229880 119100 230120 119120
rect 230380 119100 230620 119120
rect 230880 119100 231120 119120
rect 231380 119100 232000 119120
rect 214000 118900 232000 119100
rect 214000 118880 214120 118900
rect 214380 118880 214620 118900
rect 214880 118880 215120 118900
rect 215380 118880 215620 118900
rect 215880 118880 216120 118900
rect 216380 118880 216620 118900
rect 216880 118880 217120 118900
rect 217380 118880 217620 118900
rect 217880 118880 218120 118900
rect 218380 118880 218620 118900
rect 218880 118880 219120 118900
rect 219380 118880 219620 118900
rect 219880 118880 220120 118900
rect 220380 118880 220620 118900
rect 220880 118880 221120 118900
rect 221380 118880 221620 118900
rect 221880 118880 222120 118900
rect 222380 118880 222620 118900
rect 222880 118880 223120 118900
rect 223380 118880 223620 118900
rect 223880 118880 224120 118900
rect 224380 118880 224620 118900
rect 224880 118880 225120 118900
rect 225380 118880 225620 118900
rect 225880 118880 226120 118900
rect 226380 118880 226620 118900
rect 226880 118880 227120 118900
rect 227380 118880 227620 118900
rect 227880 118880 228120 118900
rect 228380 118880 228620 118900
rect 228880 118880 229120 118900
rect 229380 118880 229620 118900
rect 229880 118880 230120 118900
rect 230380 118880 230620 118900
rect 230880 118880 231120 118900
rect 231380 118880 231620 118900
rect 231880 118880 232000 118900
rect 214000 118620 214100 118880
rect 214400 118620 214600 118880
rect 214900 118620 215100 118880
rect 215400 118620 215600 118880
rect 215900 118620 216100 118880
rect 216400 118620 216600 118880
rect 216900 118620 217100 118880
rect 217400 118620 217600 118880
rect 217900 118620 218100 118880
rect 218400 118620 218600 118880
rect 218900 118620 219100 118880
rect 219400 118620 219600 118880
rect 219900 118620 220100 118880
rect 220400 118620 220600 118880
rect 220900 118620 221100 118880
rect 221400 118620 221600 118880
rect 221900 118620 222100 118880
rect 222400 118620 222600 118880
rect 222900 118620 223100 118880
rect 223400 118620 223600 118880
rect 223900 118620 224100 118880
rect 224400 118620 224600 118880
rect 224900 118620 225100 118880
rect 225400 118620 225600 118880
rect 225900 118620 226100 118880
rect 226400 118620 226600 118880
rect 226900 118620 227100 118880
rect 227400 118620 227600 118880
rect 227900 118620 228100 118880
rect 228400 118620 228600 118880
rect 228900 118620 229100 118880
rect 229400 118620 229600 118880
rect 229900 118620 230100 118880
rect 230400 118620 230600 118880
rect 230900 118620 231100 118880
rect 231400 118620 231600 118880
rect 231900 118620 232000 118880
rect 214000 118600 214120 118620
rect 214380 118600 214620 118620
rect 214880 118600 215120 118620
rect 215380 118600 215620 118620
rect 215880 118600 216120 118620
rect 216380 118600 216620 118620
rect 216880 118600 217120 118620
rect 217380 118600 217620 118620
rect 217880 118600 218120 118620
rect 218380 118600 218620 118620
rect 218880 118600 219120 118620
rect 219380 118600 219620 118620
rect 219880 118600 220120 118620
rect 220380 118600 220620 118620
rect 220880 118600 221120 118620
rect 221380 118600 221620 118620
rect 221880 118600 222120 118620
rect 222380 118600 222620 118620
rect 222880 118600 223120 118620
rect 223380 118600 223620 118620
rect 223880 118600 224120 118620
rect 224380 118600 224620 118620
rect 224880 118600 225120 118620
rect 225380 118600 225620 118620
rect 225880 118600 226120 118620
rect 226380 118600 226620 118620
rect 226880 118600 227120 118620
rect 227380 118600 227620 118620
rect 227880 118600 228120 118620
rect 228380 118600 228620 118620
rect 228880 118600 229120 118620
rect 229380 118600 229620 118620
rect 229880 118600 230120 118620
rect 230380 118600 230620 118620
rect 230880 118600 231120 118620
rect 231380 118600 231620 118620
rect 231880 118600 232000 118620
rect 214000 118400 232000 118600
rect 214000 118380 214120 118400
rect 214380 118380 214620 118400
rect 214880 118380 215120 118400
rect 215380 118380 215620 118400
rect 215880 118380 216120 118400
rect 216380 118380 216620 118400
rect 216880 118380 217120 118400
rect 217380 118380 217620 118400
rect 217880 118380 218120 118400
rect 218380 118380 218620 118400
rect 218880 118380 219120 118400
rect 219380 118380 219620 118400
rect 219880 118380 220120 118400
rect 220380 118380 220620 118400
rect 220880 118380 221120 118400
rect 221380 118380 221620 118400
rect 221880 118380 222120 118400
rect 222380 118380 222620 118400
rect 222880 118380 223120 118400
rect 223380 118380 223620 118400
rect 223880 118380 224120 118400
rect 224380 118380 224620 118400
rect 224880 118380 225120 118400
rect 225380 118380 225620 118400
rect 225880 118380 226120 118400
rect 226380 118380 226620 118400
rect 226880 118380 227120 118400
rect 227380 118380 227620 118400
rect 227880 118380 228120 118400
rect 228380 118380 228620 118400
rect 228880 118380 229120 118400
rect 229380 118380 229620 118400
rect 229880 118380 230120 118400
rect 230380 118380 230620 118400
rect 230880 118380 231120 118400
rect 231380 118380 231620 118400
rect 231880 118380 232000 118400
rect 214000 118120 214100 118380
rect 214400 118120 214600 118380
rect 214900 118120 215100 118380
rect 215400 118120 215600 118380
rect 215900 118120 216100 118380
rect 216400 118120 216600 118380
rect 216900 118120 217100 118380
rect 217400 118120 217600 118380
rect 217900 118120 218100 118380
rect 218400 118120 218600 118380
rect 218900 118120 219100 118380
rect 219400 118120 219600 118380
rect 219900 118120 220100 118380
rect 220400 118120 220600 118380
rect 220900 118120 221100 118380
rect 221400 118120 221600 118380
rect 221900 118120 222100 118380
rect 222400 118120 222600 118380
rect 222900 118120 223100 118380
rect 223400 118120 223600 118380
rect 223900 118120 224100 118380
rect 224400 118120 224600 118380
rect 224900 118120 225100 118380
rect 225400 118120 225600 118380
rect 225900 118120 226100 118380
rect 226400 118120 226600 118380
rect 226900 118120 227100 118380
rect 227400 118120 227600 118380
rect 227900 118120 228100 118380
rect 228400 118120 228600 118380
rect 228900 118120 229100 118380
rect 229400 118120 229600 118380
rect 229900 118120 230100 118380
rect 230400 118120 230600 118380
rect 230900 118120 231100 118380
rect 231400 118120 231600 118380
rect 231900 118120 232000 118380
rect 214000 118100 214120 118120
rect 214380 118100 214620 118120
rect 214880 118100 215120 118120
rect 215380 118100 215620 118120
rect 215880 118100 216120 118120
rect 216380 118100 216620 118120
rect 216880 118100 217120 118120
rect 217380 118100 217620 118120
rect 217880 118100 218120 118120
rect 218380 118100 218620 118120
rect 218880 118100 219120 118120
rect 219380 118100 219620 118120
rect 219880 118100 220120 118120
rect 220380 118100 220620 118120
rect 220880 118100 221120 118120
rect 221380 118100 221620 118120
rect 221880 118100 222120 118120
rect 222380 118100 222620 118120
rect 222880 118100 223120 118120
rect 223380 118100 223620 118120
rect 223880 118100 224120 118120
rect 224380 118100 224620 118120
rect 224880 118100 225120 118120
rect 225380 118100 225620 118120
rect 225880 118100 226120 118120
rect 226380 118100 226620 118120
rect 226880 118100 227120 118120
rect 227380 118100 227620 118120
rect 227880 118100 228120 118120
rect 228380 118100 228620 118120
rect 228880 118100 229120 118120
rect 229380 118100 229620 118120
rect 229880 118100 230120 118120
rect 230380 118100 230620 118120
rect 230880 118100 231120 118120
rect 231380 118100 231620 118120
rect 231880 118100 232000 118120
rect 214000 117900 232000 118100
rect 214000 117880 214120 117900
rect 214380 117880 214620 117900
rect 214880 117880 215120 117900
rect 215380 117880 215620 117900
rect 215880 117880 216120 117900
rect 216380 117880 216620 117900
rect 216880 117880 217120 117900
rect 217380 117880 217620 117900
rect 217880 117880 218120 117900
rect 218380 117880 218620 117900
rect 218880 117880 219120 117900
rect 219380 117880 219620 117900
rect 219880 117880 220120 117900
rect 220380 117880 220620 117900
rect 220880 117880 221120 117900
rect 221380 117880 221620 117900
rect 221880 117880 222120 117900
rect 222380 117880 222620 117900
rect 222880 117880 223120 117900
rect 223380 117880 223620 117900
rect 223880 117880 224120 117900
rect 224380 117880 224620 117900
rect 224880 117880 225120 117900
rect 225380 117880 225620 117900
rect 225880 117880 226120 117900
rect 226380 117880 226620 117900
rect 226880 117880 227120 117900
rect 227380 117880 227620 117900
rect 227880 117880 228120 117900
rect 228380 117880 228620 117900
rect 228880 117880 229120 117900
rect 229380 117880 229620 117900
rect 229880 117880 230120 117900
rect 230380 117880 230620 117900
rect 230880 117880 231120 117900
rect 231380 117880 231620 117900
rect 231880 117880 232000 117900
rect 214000 117620 214100 117880
rect 214400 117620 214600 117880
rect 214900 117620 215100 117880
rect 215400 117620 215600 117880
rect 215900 117620 216100 117880
rect 216400 117620 216600 117880
rect 216900 117620 217100 117880
rect 217400 117620 217600 117880
rect 217900 117620 218100 117880
rect 218400 117620 218600 117880
rect 218900 117620 219100 117880
rect 219400 117620 219600 117880
rect 219900 117620 220100 117880
rect 220400 117620 220600 117880
rect 220900 117620 221100 117880
rect 221400 117620 221600 117880
rect 221900 117620 222100 117880
rect 222400 117620 222600 117880
rect 222900 117620 223100 117880
rect 223400 117620 223600 117880
rect 223900 117620 224100 117880
rect 224400 117620 224600 117880
rect 224900 117620 225100 117880
rect 225400 117620 225600 117880
rect 225900 117620 226100 117880
rect 226400 117620 226600 117880
rect 226900 117620 227100 117880
rect 227400 117620 227600 117880
rect 227900 117620 228100 117880
rect 228400 117620 228600 117880
rect 228900 117620 229100 117880
rect 229400 117620 229600 117880
rect 229900 117620 230100 117880
rect 230400 117620 230600 117880
rect 230900 117620 231100 117880
rect 231400 117620 231600 117880
rect 231900 117620 232000 117880
rect 214000 117600 214120 117620
rect 214380 117600 214620 117620
rect 214880 117600 215120 117620
rect 215380 117600 215620 117620
rect 215880 117600 216120 117620
rect 216380 117600 216620 117620
rect 216880 117600 217120 117620
rect 217380 117600 217620 117620
rect 217880 117600 218120 117620
rect 218380 117600 218620 117620
rect 218880 117600 219120 117620
rect 219380 117600 219620 117620
rect 219880 117600 220120 117620
rect 220380 117600 220620 117620
rect 220880 117600 221120 117620
rect 221380 117600 221620 117620
rect 221880 117600 222120 117620
rect 222380 117600 222620 117620
rect 222880 117600 223120 117620
rect 223380 117600 223620 117620
rect 223880 117600 224120 117620
rect 224380 117600 224620 117620
rect 224880 117600 225120 117620
rect 225380 117600 225620 117620
rect 225880 117600 226120 117620
rect 226380 117600 226620 117620
rect 226880 117600 227120 117620
rect 227380 117600 227620 117620
rect 227880 117600 228120 117620
rect 228380 117600 228620 117620
rect 228880 117600 229120 117620
rect 229380 117600 229620 117620
rect 229880 117600 230120 117620
rect 230380 117600 230620 117620
rect 230880 117600 231120 117620
rect 231380 117600 231620 117620
rect 231880 117600 232000 117620
rect 214000 117400 232000 117600
rect 214000 117380 214120 117400
rect 214380 117380 214620 117400
rect 214880 117380 215120 117400
rect 215380 117380 215620 117400
rect 215880 117380 216120 117400
rect 216380 117380 216620 117400
rect 216880 117380 217120 117400
rect 217380 117380 217620 117400
rect 217880 117380 218120 117400
rect 218380 117380 218620 117400
rect 218880 117380 219120 117400
rect 219380 117380 219620 117400
rect 219880 117380 220120 117400
rect 220380 117380 220620 117400
rect 220880 117380 221120 117400
rect 221380 117380 221620 117400
rect 221880 117380 222120 117400
rect 222380 117380 222620 117400
rect 222880 117380 223120 117400
rect 223380 117380 223620 117400
rect 223880 117380 224120 117400
rect 224380 117380 224620 117400
rect 224880 117380 225120 117400
rect 225380 117380 225620 117400
rect 225880 117380 226120 117400
rect 226380 117380 226620 117400
rect 226880 117380 227120 117400
rect 227380 117380 227620 117400
rect 227880 117380 228120 117400
rect 228380 117380 228620 117400
rect 228880 117380 229120 117400
rect 229380 117380 229620 117400
rect 229880 117380 230120 117400
rect 230380 117380 230620 117400
rect 230880 117380 231120 117400
rect 231380 117380 231620 117400
rect 231880 117380 232000 117400
rect 214000 117120 214100 117380
rect 214400 117120 214600 117380
rect 214900 117120 215100 117380
rect 215400 117120 215600 117380
rect 215900 117120 216100 117380
rect 216400 117120 216600 117380
rect 216900 117120 217100 117380
rect 217400 117120 217600 117380
rect 217900 117120 218100 117380
rect 218400 117120 218600 117380
rect 218900 117120 219100 117380
rect 219400 117120 219600 117380
rect 219900 117120 220100 117380
rect 220400 117120 220600 117380
rect 220900 117120 221100 117380
rect 221400 117120 221600 117380
rect 221900 117120 222100 117380
rect 222400 117120 222600 117380
rect 222900 117120 223100 117380
rect 223400 117120 223600 117380
rect 223900 117120 224100 117380
rect 224400 117120 224600 117380
rect 224900 117120 225100 117380
rect 225400 117120 225600 117380
rect 225900 117120 226100 117380
rect 226400 117120 226600 117380
rect 226900 117120 227100 117380
rect 227400 117120 227600 117380
rect 227900 117120 228100 117380
rect 228400 117120 228600 117380
rect 228900 117120 229100 117380
rect 229400 117120 229600 117380
rect 229900 117120 230100 117380
rect 230400 117120 230600 117380
rect 230900 117120 231100 117380
rect 231400 117120 231600 117380
rect 231900 117120 232000 117380
rect 214000 117100 214120 117120
rect 214380 117100 214620 117120
rect 214880 117100 215120 117120
rect 215380 117100 215620 117120
rect 215880 117100 216120 117120
rect 216380 117100 216620 117120
rect 216880 117100 217120 117120
rect 217380 117100 217620 117120
rect 217880 117100 218120 117120
rect 218380 117100 218620 117120
rect 218880 117100 219120 117120
rect 219380 117100 219620 117120
rect 219880 117100 220120 117120
rect 220380 117100 220620 117120
rect 220880 117100 221120 117120
rect 221380 117100 221620 117120
rect 221880 117100 222120 117120
rect 222380 117100 222620 117120
rect 222880 117100 223120 117120
rect 223380 117100 223620 117120
rect 223880 117100 224120 117120
rect 224380 117100 224620 117120
rect 224880 117100 225120 117120
rect 225380 117100 225620 117120
rect 225880 117100 226120 117120
rect 226380 117100 226620 117120
rect 226880 117100 227120 117120
rect 227380 117100 227620 117120
rect 227880 117100 228120 117120
rect 228380 117100 228620 117120
rect 228880 117100 229120 117120
rect 229380 117100 229620 117120
rect 229880 117100 230120 117120
rect 230380 117100 230620 117120
rect 230880 117100 231120 117120
rect 231380 117100 231620 117120
rect 231880 117100 232000 117120
rect 214000 116900 232000 117100
rect 214000 116880 214120 116900
rect 214380 116880 214620 116900
rect 214880 116880 215120 116900
rect 215380 116880 215620 116900
rect 215880 116880 216120 116900
rect 216380 116880 216620 116900
rect 216880 116880 217120 116900
rect 217380 116880 217620 116900
rect 217880 116880 218120 116900
rect 218380 116880 218620 116900
rect 218880 116880 219120 116900
rect 219380 116880 219620 116900
rect 219880 116880 220120 116900
rect 220380 116880 220620 116900
rect 220880 116880 221120 116900
rect 221380 116880 221620 116900
rect 221880 116880 222120 116900
rect 222380 116880 222620 116900
rect 222880 116880 223120 116900
rect 223380 116880 223620 116900
rect 223880 116880 224120 116900
rect 224380 116880 224620 116900
rect 224880 116880 225120 116900
rect 225380 116880 225620 116900
rect 225880 116880 226120 116900
rect 226380 116880 226620 116900
rect 226880 116880 227120 116900
rect 227380 116880 227620 116900
rect 227880 116880 228120 116900
rect 228380 116880 228620 116900
rect 228880 116880 229120 116900
rect 229380 116880 229620 116900
rect 229880 116880 230120 116900
rect 230380 116880 230620 116900
rect 230880 116880 231120 116900
rect 231380 116880 231620 116900
rect 231880 116880 232000 116900
rect 214000 116620 214100 116880
rect 214400 116620 214600 116880
rect 214900 116620 215100 116880
rect 215400 116620 215600 116880
rect 215900 116620 216100 116880
rect 216400 116620 216600 116880
rect 216900 116620 217100 116880
rect 217400 116620 217600 116880
rect 217900 116620 218100 116880
rect 218400 116620 218600 116880
rect 218900 116620 219100 116880
rect 219400 116620 219600 116880
rect 219900 116620 220100 116880
rect 220400 116620 220600 116880
rect 220900 116620 221100 116880
rect 221400 116620 221600 116880
rect 221900 116620 222100 116880
rect 222400 116620 222600 116880
rect 222900 116620 223100 116880
rect 223400 116620 223600 116880
rect 223900 116620 224100 116880
rect 224400 116620 224600 116880
rect 224900 116620 225100 116880
rect 225400 116620 225600 116880
rect 225900 116620 226100 116880
rect 226400 116620 226600 116880
rect 226900 116620 227100 116880
rect 227400 116620 227600 116880
rect 227900 116620 228100 116880
rect 228400 116620 228600 116880
rect 228900 116620 229100 116880
rect 229400 116620 229600 116880
rect 229900 116620 230100 116880
rect 230400 116620 230600 116880
rect 230900 116620 231100 116880
rect 231400 116620 231600 116880
rect 231900 116620 232000 116880
rect 214000 116600 214120 116620
rect 214380 116600 214620 116620
rect 214880 116600 215120 116620
rect 215380 116600 215620 116620
rect 215880 116600 216120 116620
rect 216380 116600 216620 116620
rect 216880 116600 217120 116620
rect 217380 116600 217620 116620
rect 217880 116600 218120 116620
rect 218380 116600 218620 116620
rect 218880 116600 219120 116620
rect 219380 116600 219620 116620
rect 219880 116600 220120 116620
rect 220380 116600 220620 116620
rect 220880 116600 221120 116620
rect 221380 116600 221620 116620
rect 221880 116600 222120 116620
rect 222380 116600 222620 116620
rect 222880 116600 223120 116620
rect 223380 116600 223620 116620
rect 223880 116600 224120 116620
rect 224380 116600 224620 116620
rect 224880 116600 225120 116620
rect 225380 116600 225620 116620
rect 225880 116600 226120 116620
rect 226380 116600 226620 116620
rect 226880 116600 227120 116620
rect 227380 116600 227620 116620
rect 227880 116600 228120 116620
rect 228380 116600 228620 116620
rect 228880 116600 229120 116620
rect 229380 116600 229620 116620
rect 229880 116600 230120 116620
rect 230380 116600 230620 116620
rect 230880 116600 231120 116620
rect 231380 116600 231620 116620
rect 231880 116600 232000 116620
rect 214000 116400 232000 116600
rect 214000 116380 214120 116400
rect 214380 116380 214620 116400
rect 214880 116380 215120 116400
rect 215380 116380 215620 116400
rect 215880 116380 216120 116400
rect 216380 116380 216620 116400
rect 216880 116380 217120 116400
rect 217380 116380 217620 116400
rect 217880 116380 218120 116400
rect 218380 116380 218620 116400
rect 218880 116380 219120 116400
rect 219380 116380 219620 116400
rect 219880 116380 220120 116400
rect 220380 116380 220620 116400
rect 220880 116380 221120 116400
rect 221380 116380 221620 116400
rect 221880 116380 222120 116400
rect 222380 116380 222620 116400
rect 222880 116380 223120 116400
rect 223380 116380 223620 116400
rect 223880 116380 224120 116400
rect 224380 116380 224620 116400
rect 224880 116380 225120 116400
rect 225380 116380 225620 116400
rect 225880 116380 226120 116400
rect 226380 116380 226620 116400
rect 226880 116380 227120 116400
rect 227380 116380 227620 116400
rect 227880 116380 228120 116400
rect 228380 116380 228620 116400
rect 228880 116380 229120 116400
rect 229380 116380 229620 116400
rect 229880 116380 230120 116400
rect 230380 116380 230620 116400
rect 230880 116380 231120 116400
rect 231380 116380 231620 116400
rect 231880 116380 232000 116400
rect 214000 116120 214100 116380
rect 214400 116120 214600 116380
rect 214900 116120 215100 116380
rect 215400 116120 215600 116380
rect 215900 116120 216100 116380
rect 216400 116120 216600 116380
rect 216900 116120 217100 116380
rect 217400 116120 217600 116380
rect 217900 116120 218100 116380
rect 218400 116120 218600 116380
rect 218900 116120 219100 116380
rect 219400 116120 219600 116380
rect 219900 116120 220100 116380
rect 220400 116120 220600 116380
rect 220900 116120 221100 116380
rect 221400 116120 221600 116380
rect 221900 116120 222100 116380
rect 222400 116120 222600 116380
rect 222900 116120 223100 116380
rect 223400 116120 223600 116380
rect 223900 116120 224100 116380
rect 224400 116120 224600 116380
rect 224900 116120 225100 116380
rect 225400 116120 225600 116380
rect 225900 116120 226100 116380
rect 226400 116120 226600 116380
rect 226900 116120 227100 116380
rect 227400 116120 227600 116380
rect 227900 116120 228100 116380
rect 228400 116120 228600 116380
rect 228900 116120 229100 116380
rect 229400 116120 229600 116380
rect 229900 116120 230100 116380
rect 230400 116120 230600 116380
rect 230900 116120 231100 116380
rect 231400 116120 231600 116380
rect 231900 116120 232000 116380
rect 214000 116100 214120 116120
rect 214380 116100 214620 116120
rect 214880 116100 215120 116120
rect 215380 116100 215620 116120
rect 215880 116100 216120 116120
rect 216380 116100 216620 116120
rect 216880 116100 217120 116120
rect 217380 116100 217620 116120
rect 217880 116100 218120 116120
rect 218380 116100 218620 116120
rect 218880 116100 219120 116120
rect 219380 116100 219620 116120
rect 219880 116100 220120 116120
rect 220380 116100 220620 116120
rect 220880 116100 221120 116120
rect 221380 116100 221620 116120
rect 221880 116100 222120 116120
rect 222380 116100 222620 116120
rect 222880 116100 223120 116120
rect 223380 116100 223620 116120
rect 223880 116100 224120 116120
rect 224380 116100 224620 116120
rect 224880 116100 225120 116120
rect 225380 116100 225620 116120
rect 225880 116100 226120 116120
rect 226380 116100 226620 116120
rect 226880 116100 227120 116120
rect 227380 116100 227620 116120
rect 227880 116100 228120 116120
rect 228380 116100 228620 116120
rect 228880 116100 229120 116120
rect 229380 116100 229620 116120
rect 229880 116100 230120 116120
rect 230380 116100 230620 116120
rect 230880 116100 231120 116120
rect 231380 116100 231620 116120
rect 231880 116100 232000 116120
rect 214000 115900 232000 116100
rect 214000 115880 214120 115900
rect 214380 115880 214620 115900
rect 214880 115880 215120 115900
rect 215380 115880 215620 115900
rect 215880 115880 216120 115900
rect 216380 115880 216620 115900
rect 216880 115880 217120 115900
rect 217380 115880 217620 115900
rect 217880 115880 218120 115900
rect 218380 115880 218620 115900
rect 218880 115880 219120 115900
rect 219380 115880 219620 115900
rect 219880 115880 220120 115900
rect 220380 115880 220620 115900
rect 220880 115880 221120 115900
rect 221380 115880 221620 115900
rect 221880 115880 222120 115900
rect 222380 115880 222620 115900
rect 222880 115880 223120 115900
rect 223380 115880 223620 115900
rect 223880 115880 224120 115900
rect 224380 115880 224620 115900
rect 224880 115880 225120 115900
rect 225380 115880 225620 115900
rect 225880 115880 226120 115900
rect 226380 115880 226620 115900
rect 226880 115880 227120 115900
rect 227380 115880 227620 115900
rect 227880 115880 228120 115900
rect 228380 115880 228620 115900
rect 228880 115880 229120 115900
rect 229380 115880 229620 115900
rect 229880 115880 230120 115900
rect 230380 115880 230620 115900
rect 230880 115880 231120 115900
rect 231380 115880 231620 115900
rect 231880 115880 232000 115900
rect 214000 115620 214100 115880
rect 214400 115620 214600 115880
rect 214900 115620 215100 115880
rect 215400 115620 215600 115880
rect 215900 115620 216100 115880
rect 216400 115620 216600 115880
rect 216900 115620 217100 115880
rect 217400 115620 217600 115880
rect 217900 115620 218100 115880
rect 218400 115620 218600 115880
rect 218900 115620 219100 115880
rect 219400 115620 219600 115880
rect 219900 115620 220100 115880
rect 220400 115620 220600 115880
rect 220900 115620 221100 115880
rect 221400 115620 221600 115880
rect 221900 115620 222100 115880
rect 222400 115620 222600 115880
rect 222900 115620 223100 115880
rect 223400 115620 223600 115880
rect 223900 115620 224100 115880
rect 224400 115620 224600 115880
rect 224900 115620 225100 115880
rect 225400 115620 225600 115880
rect 225900 115620 226100 115880
rect 226400 115620 226600 115880
rect 226900 115620 227100 115880
rect 227400 115620 227600 115880
rect 227900 115620 228100 115880
rect 228400 115620 228600 115880
rect 228900 115620 229100 115880
rect 229400 115620 229600 115880
rect 229900 115620 230100 115880
rect 230400 115620 230600 115880
rect 230900 115620 231100 115880
rect 231400 115620 231600 115880
rect 231900 115620 232000 115880
rect 214000 115600 214120 115620
rect 214380 115600 214620 115620
rect 214880 115600 215120 115620
rect 215380 115600 215620 115620
rect 215880 115600 216120 115620
rect 216380 115600 216620 115620
rect 216880 115600 217120 115620
rect 217380 115600 217620 115620
rect 217880 115600 218120 115620
rect 218380 115600 218620 115620
rect 218880 115600 219120 115620
rect 219380 115600 219620 115620
rect 219880 115600 220120 115620
rect 220380 115600 220620 115620
rect 220880 115600 221120 115620
rect 221380 115600 221620 115620
rect 221880 115600 222120 115620
rect 222380 115600 222620 115620
rect 222880 115600 223120 115620
rect 223380 115600 223620 115620
rect 223880 115600 224120 115620
rect 224380 115600 224620 115620
rect 224880 115600 225120 115620
rect 225380 115600 225620 115620
rect 225880 115600 226120 115620
rect 226380 115600 226620 115620
rect 226880 115600 227120 115620
rect 227380 115600 227620 115620
rect 227880 115600 228120 115620
rect 228380 115600 228620 115620
rect 228880 115600 229120 115620
rect 229380 115600 229620 115620
rect 229880 115600 230120 115620
rect 230380 115600 230620 115620
rect 230880 115600 231120 115620
rect 231380 115600 231620 115620
rect 231880 115600 232000 115620
rect 214000 115400 232000 115600
rect 214000 115380 214120 115400
rect 214380 115380 214620 115400
rect 214880 115380 215120 115400
rect 215380 115380 215620 115400
rect 215880 115380 216120 115400
rect 216380 115380 216620 115400
rect 216880 115380 217120 115400
rect 217380 115380 217620 115400
rect 217880 115380 218120 115400
rect 218380 115380 218620 115400
rect 218880 115380 219120 115400
rect 219380 115380 219620 115400
rect 219880 115380 220120 115400
rect 220380 115380 220620 115400
rect 220880 115380 221120 115400
rect 221380 115380 221620 115400
rect 221880 115380 222120 115400
rect 222380 115380 222620 115400
rect 222880 115380 223120 115400
rect 223380 115380 223620 115400
rect 223880 115380 224120 115400
rect 224380 115380 224620 115400
rect 224880 115380 225120 115400
rect 225380 115380 225620 115400
rect 225880 115380 226120 115400
rect 226380 115380 226620 115400
rect 226880 115380 227120 115400
rect 227380 115380 227620 115400
rect 227880 115380 228120 115400
rect 228380 115380 228620 115400
rect 228880 115380 229120 115400
rect 229380 115380 229620 115400
rect 229880 115380 230120 115400
rect 230380 115380 230620 115400
rect 230880 115380 231120 115400
rect 231380 115380 231620 115400
rect 231880 115380 232000 115400
rect 214000 115120 214100 115380
rect 214400 115120 214600 115380
rect 214900 115120 215100 115380
rect 215400 115120 215600 115380
rect 215900 115120 216100 115380
rect 216400 115120 216600 115380
rect 216900 115120 217100 115380
rect 217400 115120 217600 115380
rect 217900 115120 218100 115380
rect 218400 115120 218600 115380
rect 218900 115120 219100 115380
rect 219400 115120 219600 115380
rect 219900 115120 220100 115380
rect 220400 115120 220600 115380
rect 220900 115120 221100 115380
rect 221400 115120 221600 115380
rect 221900 115120 222100 115380
rect 222400 115120 222600 115380
rect 222900 115120 223100 115380
rect 223400 115120 223600 115380
rect 223900 115120 224100 115380
rect 224400 115120 224600 115380
rect 224900 115120 225100 115380
rect 225400 115120 225600 115380
rect 225900 115120 226100 115380
rect 226400 115120 226600 115380
rect 226900 115120 227100 115380
rect 227400 115120 227600 115380
rect 227900 115120 228100 115380
rect 228400 115120 228600 115380
rect 228900 115120 229100 115380
rect 229400 115120 229600 115380
rect 229900 115120 230100 115380
rect 230400 115120 230600 115380
rect 230900 115120 231100 115380
rect 231400 115120 231600 115380
rect 231900 115120 232000 115380
rect 214000 115100 214120 115120
rect 214380 115100 214620 115120
rect 214880 115100 215120 115120
rect 215380 115100 215620 115120
rect 215880 115100 216120 115120
rect 216380 115100 216620 115120
rect 216880 115100 217120 115120
rect 217380 115100 217620 115120
rect 217880 115100 218120 115120
rect 218380 115100 218620 115120
rect 218880 115100 219120 115120
rect 219380 115100 219620 115120
rect 219880 115100 220120 115120
rect 220380 115100 220620 115120
rect 220880 115100 221120 115120
rect 221380 115100 221620 115120
rect 221880 115100 222120 115120
rect 222380 115100 222620 115120
rect 222880 115100 223120 115120
rect 223380 115100 223620 115120
rect 223880 115100 224120 115120
rect 224380 115100 224620 115120
rect 224880 115100 225120 115120
rect 225380 115100 225620 115120
rect 225880 115100 226120 115120
rect 226380 115100 226620 115120
rect 226880 115100 227120 115120
rect 227380 115100 227620 115120
rect 227880 115100 228120 115120
rect 228380 115100 228620 115120
rect 228880 115100 229120 115120
rect 229380 115100 229620 115120
rect 229880 115100 230120 115120
rect 230380 115100 230620 115120
rect 230880 115100 231120 115120
rect 231380 115100 231620 115120
rect 231880 115100 232000 115120
rect 214000 114900 232000 115100
rect 214000 114880 214120 114900
rect 214380 114880 214620 114900
rect 214880 114880 215120 114900
rect 215380 114880 215620 114900
rect 215880 114880 216120 114900
rect 216380 114880 216620 114900
rect 216880 114880 217120 114900
rect 217380 114880 217620 114900
rect 217880 114880 218120 114900
rect 218380 114880 218620 114900
rect 218880 114880 219120 114900
rect 219380 114880 219620 114900
rect 219880 114880 220120 114900
rect 220380 114880 220620 114900
rect 220880 114880 221120 114900
rect 221380 114880 221620 114900
rect 221880 114880 222120 114900
rect 222380 114880 222620 114900
rect 222880 114880 223120 114900
rect 223380 114880 223620 114900
rect 223880 114880 224120 114900
rect 224380 114880 224620 114900
rect 224880 114880 225120 114900
rect 225380 114880 225620 114900
rect 225880 114880 226120 114900
rect 226380 114880 226620 114900
rect 226880 114880 227120 114900
rect 227380 114880 227620 114900
rect 227880 114880 228120 114900
rect 228380 114880 228620 114900
rect 228880 114880 229120 114900
rect 229380 114880 229620 114900
rect 229880 114880 230120 114900
rect 230380 114880 230620 114900
rect 230880 114880 231120 114900
rect 231380 114880 231620 114900
rect 231880 114880 232000 114900
rect 214000 114620 214100 114880
rect 214400 114620 214600 114880
rect 214900 114620 215100 114880
rect 215400 114620 215600 114880
rect 215900 114620 216100 114880
rect 216400 114620 216600 114880
rect 216900 114620 217100 114880
rect 217400 114620 217600 114880
rect 217900 114620 218100 114880
rect 218400 114620 218600 114880
rect 218900 114620 219100 114880
rect 219400 114620 219600 114880
rect 219900 114620 220100 114880
rect 220400 114620 220600 114880
rect 220900 114620 221100 114880
rect 221400 114620 221600 114880
rect 221900 114620 222100 114880
rect 222400 114620 222600 114880
rect 222900 114620 223100 114880
rect 223400 114620 223600 114880
rect 223900 114620 224100 114880
rect 224400 114620 224600 114880
rect 224900 114620 225100 114880
rect 225400 114620 225600 114880
rect 225900 114620 226100 114880
rect 226400 114620 226600 114880
rect 226900 114620 227100 114880
rect 227400 114620 227600 114880
rect 227900 114620 228100 114880
rect 228400 114620 228600 114880
rect 228900 114620 229100 114880
rect 229400 114620 229600 114880
rect 229900 114620 230100 114880
rect 230400 114620 230600 114880
rect 230900 114620 231100 114880
rect 231400 114620 231600 114880
rect 231900 114620 232000 114880
rect 214000 114600 214120 114620
rect 214380 114600 214620 114620
rect 214880 114600 215120 114620
rect 215380 114600 215620 114620
rect 215880 114600 216120 114620
rect 216380 114600 216620 114620
rect 216880 114600 217120 114620
rect 217380 114600 217620 114620
rect 217880 114600 218120 114620
rect 218380 114600 218620 114620
rect 218880 114600 219120 114620
rect 219380 114600 219620 114620
rect 219880 114600 220120 114620
rect 220380 114600 220620 114620
rect 220880 114600 221120 114620
rect 221380 114600 221620 114620
rect 221880 114600 222120 114620
rect 222380 114600 222620 114620
rect 222880 114600 223120 114620
rect 223380 114600 223620 114620
rect 223880 114600 224120 114620
rect 224380 114600 224620 114620
rect 224880 114600 225120 114620
rect 225380 114600 225620 114620
rect 225880 114600 226120 114620
rect 226380 114600 226620 114620
rect 226880 114600 227120 114620
rect 227380 114600 227620 114620
rect 227880 114600 228120 114620
rect 228380 114600 228620 114620
rect 228880 114600 229120 114620
rect 229380 114600 229620 114620
rect 229880 114600 230120 114620
rect 230380 114600 230620 114620
rect 230880 114600 231120 114620
rect 231380 114600 231620 114620
rect 231880 114600 232000 114620
rect 214000 114400 232000 114600
rect 214000 114380 214120 114400
rect 214380 114380 214620 114400
rect 214880 114380 215120 114400
rect 215380 114380 215620 114400
rect 215880 114380 216120 114400
rect 216380 114380 216620 114400
rect 216880 114380 217120 114400
rect 217380 114380 217620 114400
rect 217880 114380 218120 114400
rect 218380 114380 218620 114400
rect 218880 114380 219120 114400
rect 219380 114380 219620 114400
rect 219880 114380 220120 114400
rect 220380 114380 220620 114400
rect 220880 114380 221120 114400
rect 221380 114380 221620 114400
rect 221880 114380 222120 114400
rect 222380 114380 222620 114400
rect 222880 114380 223120 114400
rect 223380 114380 223620 114400
rect 223880 114380 224120 114400
rect 224380 114380 224620 114400
rect 224880 114380 225120 114400
rect 225380 114380 225620 114400
rect 225880 114380 226120 114400
rect 226380 114380 226620 114400
rect 226880 114380 227120 114400
rect 227380 114380 227620 114400
rect 227880 114380 228120 114400
rect 228380 114380 228620 114400
rect 228880 114380 229120 114400
rect 229380 114380 229620 114400
rect 229880 114380 230120 114400
rect 230380 114380 230620 114400
rect 230880 114380 231120 114400
rect 231380 114380 231620 114400
rect 231880 114380 232000 114400
rect 214000 114120 214100 114380
rect 214400 114120 214600 114380
rect 214900 114120 215100 114380
rect 215400 114120 215600 114380
rect 215900 114120 216100 114380
rect 216400 114120 216600 114380
rect 216900 114120 217100 114380
rect 217400 114120 217600 114380
rect 217900 114120 218100 114380
rect 218400 114120 218600 114380
rect 218900 114120 219100 114380
rect 219400 114120 219600 114380
rect 219900 114120 220100 114380
rect 220400 114120 220600 114380
rect 220900 114120 221100 114380
rect 221400 114120 221600 114380
rect 221900 114120 222100 114380
rect 222400 114120 222600 114380
rect 222900 114120 223100 114380
rect 223400 114120 223600 114380
rect 223900 114120 224100 114380
rect 224400 114120 224600 114380
rect 224900 114120 225100 114380
rect 225400 114120 225600 114380
rect 225900 114120 226100 114380
rect 226400 114120 226600 114380
rect 226900 114120 227100 114380
rect 227400 114120 227600 114380
rect 227900 114120 228100 114380
rect 228400 114120 228600 114380
rect 228900 114120 229100 114380
rect 229400 114120 229600 114380
rect 229900 114120 230100 114380
rect 230400 114120 230600 114380
rect 230900 114120 231100 114380
rect 231400 114120 231600 114380
rect 231900 114120 232000 114380
rect 214000 114100 214120 114120
rect 214380 114100 214620 114120
rect 214880 114100 215120 114120
rect 215380 114100 215620 114120
rect 215880 114100 216120 114120
rect 216380 114100 216620 114120
rect 216880 114100 217120 114120
rect 217380 114100 217620 114120
rect 217880 114100 218120 114120
rect 218380 114100 218620 114120
rect 218880 114100 219120 114120
rect 219380 114100 219620 114120
rect 219880 114100 220120 114120
rect 220380 114100 220620 114120
rect 220880 114100 221120 114120
rect 221380 114100 221620 114120
rect 221880 114100 222120 114120
rect 222380 114100 222620 114120
rect 222880 114100 223120 114120
rect 223380 114100 223620 114120
rect 223880 114100 224120 114120
rect 224380 114100 224620 114120
rect 224880 114100 225120 114120
rect 225380 114100 225620 114120
rect 225880 114100 226120 114120
rect 226380 114100 226620 114120
rect 226880 114100 227120 114120
rect 227380 114100 227620 114120
rect 227880 114100 228120 114120
rect 228380 114100 228620 114120
rect 228880 114100 229120 114120
rect 229380 114100 229620 114120
rect 229880 114100 230120 114120
rect 230380 114100 230620 114120
rect 230880 114100 231120 114120
rect 231380 114100 231620 114120
rect 231880 114100 232000 114120
rect 214000 114000 232000 114100
rect 178000 113900 232000 114000
rect 178000 113880 178120 113900
rect 178380 113880 178620 113900
rect 178880 113880 179120 113900
rect 179380 113880 179620 113900
rect 179880 113880 180120 113900
rect 180380 113880 180620 113900
rect 180880 113880 181120 113900
rect 181380 113880 181620 113900
rect 181880 113880 182120 113900
rect 182380 113880 182620 113900
rect 182880 113880 183120 113900
rect 183380 113880 183620 113900
rect 183880 113880 184120 113900
rect 184380 113880 184620 113900
rect 184880 113880 185120 113900
rect 185380 113880 185620 113900
rect 185880 113880 186120 113900
rect 186380 113880 186620 113900
rect 186880 113880 187120 113900
rect 187380 113880 187620 113900
rect 187880 113880 188120 113900
rect 188380 113880 188620 113900
rect 188880 113880 189120 113900
rect 189380 113880 189620 113900
rect 189880 113880 190120 113900
rect 190380 113880 190620 113900
rect 190880 113880 191120 113900
rect 191380 113880 191620 113900
rect 191880 113880 192120 113900
rect 192380 113880 192620 113900
rect 192880 113880 193120 113900
rect 193380 113880 193620 113900
rect 193880 113880 194120 113900
rect 194380 113880 194620 113900
rect 194880 113880 195120 113900
rect 195380 113880 195620 113900
rect 195880 113880 196120 113900
rect 196380 113880 196620 113900
rect 196880 113880 197120 113900
rect 197380 113880 197620 113900
rect 197880 113880 198120 113900
rect 198380 113880 198620 113900
rect 198880 113880 199120 113900
rect 199380 113880 199620 113900
rect 199880 113880 200120 113900
rect 200380 113880 200620 113900
rect 200880 113880 201120 113900
rect 201380 113880 201620 113900
rect 201880 113880 202120 113900
rect 202380 113880 202620 113900
rect 202880 113880 203120 113900
rect 203380 113880 203620 113900
rect 203880 113880 204120 113900
rect 204380 113880 204620 113900
rect 204880 113880 205120 113900
rect 205380 113880 205620 113900
rect 205880 113880 206120 113900
rect 206380 113880 206620 113900
rect 206880 113880 207120 113900
rect 207380 113880 207620 113900
rect 207880 113880 208120 113900
rect 208380 113880 208620 113900
rect 208880 113880 209120 113900
rect 209380 113880 209620 113900
rect 209880 113880 210120 113900
rect 210380 113880 210620 113900
rect 210880 113880 211120 113900
rect 211380 113880 211620 113900
rect 211880 113880 212120 113900
rect 212380 113880 212620 113900
rect 212880 113880 213120 113900
rect 213380 113880 213620 113900
rect 213880 113880 214120 113900
rect 214380 113880 214620 113900
rect 214880 113880 215120 113900
rect 215380 113880 215620 113900
rect 215880 113880 216120 113900
rect 216380 113880 216620 113900
rect 216880 113880 217120 113900
rect 217380 113880 217620 113900
rect 217880 113880 218120 113900
rect 218380 113880 218620 113900
rect 218880 113880 219120 113900
rect 219380 113880 219620 113900
rect 219880 113880 220120 113900
rect 220380 113880 220620 113900
rect 220880 113880 221120 113900
rect 221380 113880 221620 113900
rect 221880 113880 222120 113900
rect 222380 113880 222620 113900
rect 222880 113880 223120 113900
rect 223380 113880 223620 113900
rect 223880 113880 224120 113900
rect 224380 113880 224620 113900
rect 224880 113880 225120 113900
rect 225380 113880 225620 113900
rect 225880 113880 226120 113900
rect 226380 113880 226620 113900
rect 226880 113880 227120 113900
rect 227380 113880 227620 113900
rect 227880 113880 228120 113900
rect 228380 113880 228620 113900
rect 228880 113880 229120 113900
rect 229380 113880 229620 113900
rect 229880 113880 230120 113900
rect 230380 113880 230620 113900
rect 230880 113880 231120 113900
rect 231380 113880 231620 113900
rect 231880 113880 232000 113900
rect 178000 113620 178100 113880
rect 178400 113620 178600 113880
rect 178900 113620 179100 113880
rect 179400 113620 179600 113880
rect 179900 113620 180100 113880
rect 180400 113620 180600 113880
rect 180900 113620 181100 113880
rect 181400 113620 181600 113880
rect 181900 113620 182100 113880
rect 182400 113620 182600 113880
rect 182900 113620 183100 113880
rect 183400 113620 183600 113880
rect 183900 113620 184100 113880
rect 184400 113620 184600 113880
rect 184900 113620 185100 113880
rect 185400 113620 185600 113880
rect 185900 113620 186100 113880
rect 186400 113620 186600 113880
rect 186900 113620 187100 113880
rect 187400 113620 187600 113880
rect 187900 113620 188100 113880
rect 188400 113620 188600 113880
rect 188900 113620 189100 113880
rect 189400 113620 189600 113880
rect 189900 113620 190100 113880
rect 190400 113620 190600 113880
rect 190900 113620 191100 113880
rect 191400 113620 191600 113880
rect 191900 113620 192100 113880
rect 192400 113620 192600 113880
rect 192900 113620 193100 113880
rect 193400 113620 193600 113880
rect 193900 113620 194100 113880
rect 194400 113620 194600 113880
rect 194900 113620 195100 113880
rect 195400 113620 195600 113880
rect 195900 113620 196100 113880
rect 196400 113620 196600 113880
rect 196900 113620 197100 113880
rect 197400 113620 197600 113880
rect 197900 113620 198100 113880
rect 198400 113620 198600 113880
rect 198900 113620 199100 113880
rect 199400 113620 199600 113880
rect 199900 113620 200100 113880
rect 200400 113620 200600 113880
rect 200900 113620 201100 113880
rect 201400 113620 201600 113880
rect 201900 113620 202100 113880
rect 202400 113620 202600 113880
rect 202900 113620 203100 113880
rect 203400 113620 203600 113880
rect 203900 113620 204100 113880
rect 204400 113620 204600 113880
rect 204900 113620 205100 113880
rect 205400 113620 205600 113880
rect 205900 113620 206100 113880
rect 206400 113620 206600 113880
rect 206900 113620 207100 113880
rect 207400 113620 207600 113880
rect 207900 113620 208100 113880
rect 208400 113620 208600 113880
rect 208900 113620 209100 113880
rect 209400 113620 209600 113880
rect 209900 113620 210100 113880
rect 210400 113620 210600 113880
rect 210900 113620 211100 113880
rect 211400 113620 211600 113880
rect 211900 113620 212100 113880
rect 212400 113620 212600 113880
rect 212900 113620 213100 113880
rect 213400 113620 213600 113880
rect 213900 113620 214100 113880
rect 214400 113620 214600 113880
rect 214900 113620 215100 113880
rect 215400 113620 215600 113880
rect 215900 113620 216100 113880
rect 216400 113620 216600 113880
rect 216900 113620 217100 113880
rect 217400 113620 217600 113880
rect 217900 113620 218100 113880
rect 218400 113620 218600 113880
rect 218900 113620 219100 113880
rect 219400 113620 219600 113880
rect 219900 113620 220100 113880
rect 220400 113620 220600 113880
rect 220900 113620 221100 113880
rect 221400 113620 221600 113880
rect 221900 113620 222100 113880
rect 222400 113620 222600 113880
rect 222900 113620 223100 113880
rect 223400 113620 223600 113880
rect 223900 113620 224100 113880
rect 224400 113620 224600 113880
rect 224900 113620 225100 113880
rect 225400 113620 225600 113880
rect 225900 113620 226100 113880
rect 226400 113620 226600 113880
rect 226900 113620 227100 113880
rect 227400 113620 227600 113880
rect 227900 113620 228100 113880
rect 228400 113620 228600 113880
rect 228900 113620 229100 113880
rect 229400 113620 229600 113880
rect 229900 113620 230100 113880
rect 230400 113620 230600 113880
rect 230900 113620 231100 113880
rect 231400 113620 231600 113880
rect 231900 113620 232000 113880
rect 178000 113600 178120 113620
rect 178380 113600 178620 113620
rect 178880 113600 179120 113620
rect 179380 113600 179620 113620
rect 179880 113600 180120 113620
rect 180380 113600 180620 113620
rect 180880 113600 181120 113620
rect 181380 113600 181620 113620
rect 181880 113600 182120 113620
rect 182380 113600 182620 113620
rect 182880 113600 183120 113620
rect 183380 113600 183620 113620
rect 183880 113600 184120 113620
rect 184380 113600 184620 113620
rect 184880 113600 185120 113620
rect 185380 113600 185620 113620
rect 185880 113600 186120 113620
rect 186380 113600 186620 113620
rect 186880 113600 187120 113620
rect 187380 113600 187620 113620
rect 187880 113600 188120 113620
rect 188380 113600 188620 113620
rect 188880 113600 189120 113620
rect 189380 113600 189620 113620
rect 189880 113600 190120 113620
rect 190380 113600 190620 113620
rect 190880 113600 191120 113620
rect 191380 113600 191620 113620
rect 191880 113600 192120 113620
rect 192380 113600 192620 113620
rect 192880 113600 193120 113620
rect 193380 113600 193620 113620
rect 193880 113600 194120 113620
rect 194380 113600 194620 113620
rect 194880 113600 195120 113620
rect 195380 113600 195620 113620
rect 195880 113600 196120 113620
rect 196380 113600 196620 113620
rect 196880 113600 197120 113620
rect 197380 113600 197620 113620
rect 197880 113600 198120 113620
rect 198380 113600 198620 113620
rect 198880 113600 199120 113620
rect 199380 113600 199620 113620
rect 199880 113600 200120 113620
rect 200380 113600 200620 113620
rect 200880 113600 201120 113620
rect 201380 113600 201620 113620
rect 201880 113600 202120 113620
rect 202380 113600 202620 113620
rect 202880 113600 203120 113620
rect 203380 113600 203620 113620
rect 203880 113600 204120 113620
rect 204380 113600 204620 113620
rect 204880 113600 205120 113620
rect 205380 113600 205620 113620
rect 205880 113600 206120 113620
rect 206380 113600 206620 113620
rect 206880 113600 207120 113620
rect 207380 113600 207620 113620
rect 207880 113600 208120 113620
rect 208380 113600 208620 113620
rect 208880 113600 209120 113620
rect 209380 113600 209620 113620
rect 209880 113600 210120 113620
rect 210380 113600 210620 113620
rect 210880 113600 211120 113620
rect 211380 113600 211620 113620
rect 211880 113600 212120 113620
rect 212380 113600 212620 113620
rect 212880 113600 213120 113620
rect 213380 113600 213620 113620
rect 213880 113600 214120 113620
rect 214380 113600 214620 113620
rect 214880 113600 215120 113620
rect 215380 113600 215620 113620
rect 215880 113600 216120 113620
rect 216380 113600 216620 113620
rect 216880 113600 217120 113620
rect 217380 113600 217620 113620
rect 217880 113600 218120 113620
rect 218380 113600 218620 113620
rect 218880 113600 219120 113620
rect 219380 113600 219620 113620
rect 219880 113600 220120 113620
rect 220380 113600 220620 113620
rect 220880 113600 221120 113620
rect 221380 113600 221620 113620
rect 221880 113600 222120 113620
rect 222380 113600 222620 113620
rect 222880 113600 223120 113620
rect 223380 113600 223620 113620
rect 223880 113600 224120 113620
rect 224380 113600 224620 113620
rect 224880 113600 225120 113620
rect 225380 113600 225620 113620
rect 225880 113600 226120 113620
rect 226380 113600 226620 113620
rect 226880 113600 227120 113620
rect 227380 113600 227620 113620
rect 227880 113600 228120 113620
rect 228380 113600 228620 113620
rect 228880 113600 229120 113620
rect 229380 113600 229620 113620
rect 229880 113600 230120 113620
rect 230380 113600 230620 113620
rect 230880 113600 231120 113620
rect 231380 113600 231620 113620
rect 231880 113600 232000 113620
rect 178000 113400 232000 113600
rect 178000 113380 178120 113400
rect 178380 113380 178620 113400
rect 178880 113380 179120 113400
rect 179380 113380 179620 113400
rect 179880 113380 180120 113400
rect 180380 113380 180620 113400
rect 180880 113380 181120 113400
rect 181380 113380 181620 113400
rect 181880 113380 182120 113400
rect 182380 113380 182620 113400
rect 182880 113380 183120 113400
rect 183380 113380 183620 113400
rect 183880 113380 184120 113400
rect 184380 113380 184620 113400
rect 184880 113380 185120 113400
rect 185380 113380 185620 113400
rect 185880 113380 186120 113400
rect 186380 113380 186620 113400
rect 186880 113380 187120 113400
rect 187380 113380 187620 113400
rect 187880 113380 188120 113400
rect 188380 113380 188620 113400
rect 188880 113380 189120 113400
rect 189380 113380 189620 113400
rect 189880 113380 190120 113400
rect 190380 113380 190620 113400
rect 190880 113380 191120 113400
rect 191380 113380 191620 113400
rect 191880 113380 192120 113400
rect 192380 113380 192620 113400
rect 192880 113380 193120 113400
rect 193380 113380 193620 113400
rect 193880 113380 194120 113400
rect 194380 113380 194620 113400
rect 194880 113380 195120 113400
rect 195380 113380 195620 113400
rect 195880 113380 196120 113400
rect 196380 113380 196620 113400
rect 196880 113380 197120 113400
rect 197380 113380 197620 113400
rect 197880 113380 198120 113400
rect 198380 113380 198620 113400
rect 198880 113380 199120 113400
rect 199380 113380 199620 113400
rect 199880 113380 200120 113400
rect 200380 113380 200620 113400
rect 200880 113380 201120 113400
rect 201380 113380 201620 113400
rect 201880 113380 202120 113400
rect 202380 113380 202620 113400
rect 202880 113380 203120 113400
rect 203380 113380 203620 113400
rect 203880 113380 204120 113400
rect 204380 113380 204620 113400
rect 204880 113380 205120 113400
rect 205380 113380 205620 113400
rect 205880 113380 206120 113400
rect 206380 113380 206620 113400
rect 206880 113380 207120 113400
rect 207380 113380 207620 113400
rect 207880 113380 208120 113400
rect 208380 113380 208620 113400
rect 208880 113380 209120 113400
rect 209380 113380 209620 113400
rect 209880 113380 210120 113400
rect 210380 113380 210620 113400
rect 210880 113380 211120 113400
rect 211380 113380 211620 113400
rect 211880 113380 212120 113400
rect 212380 113380 212620 113400
rect 212880 113380 213120 113400
rect 213380 113380 213620 113400
rect 213880 113380 214120 113400
rect 214380 113380 214620 113400
rect 214880 113380 215120 113400
rect 215380 113380 215620 113400
rect 215880 113380 216120 113400
rect 216380 113380 216620 113400
rect 216880 113380 217120 113400
rect 217380 113380 217620 113400
rect 217880 113380 218120 113400
rect 218380 113380 218620 113400
rect 218880 113380 219120 113400
rect 219380 113380 219620 113400
rect 219880 113380 220120 113400
rect 220380 113380 220620 113400
rect 220880 113380 221120 113400
rect 221380 113380 221620 113400
rect 221880 113380 222120 113400
rect 222380 113380 222620 113400
rect 222880 113380 223120 113400
rect 223380 113380 223620 113400
rect 223880 113380 224120 113400
rect 224380 113380 224620 113400
rect 224880 113380 225120 113400
rect 225380 113380 225620 113400
rect 225880 113380 226120 113400
rect 226380 113380 226620 113400
rect 226880 113380 227120 113400
rect 227380 113380 227620 113400
rect 227880 113380 228120 113400
rect 228380 113380 228620 113400
rect 228880 113380 229120 113400
rect 229380 113380 229620 113400
rect 229880 113380 230120 113400
rect 230380 113380 230620 113400
rect 230880 113380 231120 113400
rect 231380 113380 231620 113400
rect 231880 113380 232000 113400
rect 178000 113120 178100 113380
rect 178400 113120 178600 113380
rect 178900 113120 179100 113380
rect 179400 113120 179600 113380
rect 179900 113120 180100 113380
rect 180400 113120 180600 113380
rect 180900 113120 181100 113380
rect 181400 113120 181600 113380
rect 181900 113120 182100 113380
rect 182400 113120 182600 113380
rect 182900 113120 183100 113380
rect 183400 113120 183600 113380
rect 183900 113120 184100 113380
rect 184400 113120 184600 113380
rect 184900 113120 185100 113380
rect 185400 113120 185600 113380
rect 185900 113120 186100 113380
rect 186400 113120 186600 113380
rect 186900 113120 187100 113380
rect 187400 113120 187600 113380
rect 187900 113120 188100 113380
rect 188400 113120 188600 113380
rect 188900 113120 189100 113380
rect 189400 113120 189600 113380
rect 189900 113120 190100 113380
rect 190400 113120 190600 113380
rect 190900 113120 191100 113380
rect 191400 113120 191600 113380
rect 191900 113120 192100 113380
rect 192400 113120 192600 113380
rect 192900 113120 193100 113380
rect 193400 113120 193600 113380
rect 193900 113120 194100 113380
rect 194400 113120 194600 113380
rect 194900 113120 195100 113380
rect 195400 113120 195600 113380
rect 195900 113120 196100 113380
rect 196400 113120 196600 113380
rect 196900 113120 197100 113380
rect 197400 113120 197600 113380
rect 197900 113120 198100 113380
rect 198400 113120 198600 113380
rect 198900 113120 199100 113380
rect 199400 113120 199600 113380
rect 199900 113120 200100 113380
rect 200400 113120 200600 113380
rect 200900 113120 201100 113380
rect 201400 113120 201600 113380
rect 201900 113120 202100 113380
rect 202400 113120 202600 113380
rect 202900 113120 203100 113380
rect 203400 113120 203600 113380
rect 203900 113120 204100 113380
rect 204400 113120 204600 113380
rect 204900 113120 205100 113380
rect 205400 113120 205600 113380
rect 205900 113120 206100 113380
rect 206400 113120 206600 113380
rect 206900 113120 207100 113380
rect 207400 113120 207600 113380
rect 207900 113120 208100 113380
rect 208400 113120 208600 113380
rect 208900 113120 209100 113380
rect 209400 113120 209600 113380
rect 209900 113120 210100 113380
rect 210400 113120 210600 113380
rect 210900 113120 211100 113380
rect 211400 113120 211600 113380
rect 211900 113120 212100 113380
rect 212400 113120 212600 113380
rect 212900 113120 213100 113380
rect 213400 113120 213600 113380
rect 213900 113120 214100 113380
rect 214400 113120 214600 113380
rect 214900 113120 215100 113380
rect 215400 113120 215600 113380
rect 215900 113120 216100 113380
rect 216400 113120 216600 113380
rect 216900 113120 217100 113380
rect 217400 113120 217600 113380
rect 217900 113120 218100 113380
rect 218400 113120 218600 113380
rect 218900 113120 219100 113380
rect 219400 113120 219600 113380
rect 219900 113120 220100 113380
rect 220400 113120 220600 113380
rect 220900 113120 221100 113380
rect 221400 113120 221600 113380
rect 221900 113120 222100 113380
rect 222400 113120 222600 113380
rect 222900 113120 223100 113380
rect 223400 113120 223600 113380
rect 223900 113120 224100 113380
rect 224400 113120 224600 113380
rect 224900 113120 225100 113380
rect 225400 113120 225600 113380
rect 225900 113120 226100 113380
rect 226400 113120 226600 113380
rect 226900 113120 227100 113380
rect 227400 113120 227600 113380
rect 227900 113120 228100 113380
rect 228400 113120 228600 113380
rect 228900 113120 229100 113380
rect 229400 113120 229600 113380
rect 229900 113120 230100 113380
rect 230400 113120 230600 113380
rect 230900 113120 231100 113380
rect 231400 113120 231600 113380
rect 231900 113120 232000 113380
rect 178000 113100 178120 113120
rect 178380 113100 178620 113120
rect 178880 113100 179120 113120
rect 179380 113100 179620 113120
rect 179880 113100 180120 113120
rect 180380 113100 180620 113120
rect 180880 113100 181120 113120
rect 181380 113100 181620 113120
rect 181880 113100 182120 113120
rect 182380 113100 182620 113120
rect 182880 113100 183120 113120
rect 183380 113100 183620 113120
rect 183880 113100 184120 113120
rect 184380 113100 184620 113120
rect 184880 113100 185120 113120
rect 185380 113100 185620 113120
rect 185880 113100 186120 113120
rect 186380 113100 186620 113120
rect 186880 113100 187120 113120
rect 187380 113100 187620 113120
rect 187880 113100 188120 113120
rect 188380 113100 188620 113120
rect 188880 113100 189120 113120
rect 189380 113100 189620 113120
rect 189880 113100 190120 113120
rect 190380 113100 190620 113120
rect 190880 113100 191120 113120
rect 191380 113100 191620 113120
rect 191880 113100 192120 113120
rect 192380 113100 192620 113120
rect 192880 113100 193120 113120
rect 193380 113100 193620 113120
rect 193880 113100 194120 113120
rect 194380 113100 194620 113120
rect 194880 113100 195120 113120
rect 195380 113100 195620 113120
rect 195880 113100 196120 113120
rect 196380 113100 196620 113120
rect 196880 113100 197120 113120
rect 197380 113100 197620 113120
rect 197880 113100 198120 113120
rect 198380 113100 198620 113120
rect 198880 113100 199120 113120
rect 199380 113100 199620 113120
rect 199880 113100 200120 113120
rect 200380 113100 200620 113120
rect 200880 113100 201120 113120
rect 201380 113100 201620 113120
rect 201880 113100 202120 113120
rect 202380 113100 202620 113120
rect 202880 113100 203120 113120
rect 203380 113100 203620 113120
rect 203880 113100 204120 113120
rect 204380 113100 204620 113120
rect 204880 113100 205120 113120
rect 205380 113100 205620 113120
rect 205880 113100 206120 113120
rect 206380 113100 206620 113120
rect 206880 113100 207120 113120
rect 207380 113100 207620 113120
rect 207880 113100 208120 113120
rect 208380 113100 208620 113120
rect 208880 113100 209120 113120
rect 209380 113100 209620 113120
rect 209880 113100 210120 113120
rect 210380 113100 210620 113120
rect 210880 113100 211120 113120
rect 211380 113100 211620 113120
rect 211880 113100 212120 113120
rect 212380 113100 212620 113120
rect 212880 113100 213120 113120
rect 213380 113100 213620 113120
rect 213880 113100 214120 113120
rect 214380 113100 214620 113120
rect 214880 113100 215120 113120
rect 215380 113100 215620 113120
rect 215880 113100 216120 113120
rect 216380 113100 216620 113120
rect 216880 113100 217120 113120
rect 217380 113100 217620 113120
rect 217880 113100 218120 113120
rect 218380 113100 218620 113120
rect 218880 113100 219120 113120
rect 219380 113100 219620 113120
rect 219880 113100 220120 113120
rect 220380 113100 220620 113120
rect 220880 113100 221120 113120
rect 221380 113100 221620 113120
rect 221880 113100 222120 113120
rect 222380 113100 222620 113120
rect 222880 113100 223120 113120
rect 223380 113100 223620 113120
rect 223880 113100 224120 113120
rect 224380 113100 224620 113120
rect 224880 113100 225120 113120
rect 225380 113100 225620 113120
rect 225880 113100 226120 113120
rect 226380 113100 226620 113120
rect 226880 113100 227120 113120
rect 227380 113100 227620 113120
rect 227880 113100 228120 113120
rect 228380 113100 228620 113120
rect 228880 113100 229120 113120
rect 229380 113100 229620 113120
rect 229880 113100 230120 113120
rect 230380 113100 230620 113120
rect 230880 113100 231120 113120
rect 231380 113100 231620 113120
rect 231880 113100 232000 113120
rect 178000 112900 232000 113100
rect 178000 112880 178120 112900
rect 178380 112880 178620 112900
rect 178880 112880 179120 112900
rect 179380 112880 179620 112900
rect 179880 112880 180120 112900
rect 180380 112880 180620 112900
rect 180880 112880 181120 112900
rect 181380 112880 181620 112900
rect 181880 112880 182120 112900
rect 182380 112880 182620 112900
rect 182880 112880 183120 112900
rect 183380 112880 183620 112900
rect 183880 112880 184120 112900
rect 184380 112880 184620 112900
rect 184880 112880 185120 112900
rect 185380 112880 185620 112900
rect 185880 112880 186120 112900
rect 186380 112880 186620 112900
rect 186880 112880 187120 112900
rect 187380 112880 187620 112900
rect 187880 112880 188120 112900
rect 188380 112880 188620 112900
rect 188880 112880 189120 112900
rect 189380 112880 189620 112900
rect 189880 112880 190120 112900
rect 190380 112880 190620 112900
rect 190880 112880 191120 112900
rect 191380 112880 191620 112900
rect 191880 112880 192120 112900
rect 192380 112880 192620 112900
rect 192880 112880 193120 112900
rect 193380 112880 193620 112900
rect 193880 112880 194120 112900
rect 194380 112880 194620 112900
rect 194880 112880 195120 112900
rect 195380 112880 195620 112900
rect 195880 112880 196120 112900
rect 196380 112880 196620 112900
rect 196880 112880 197120 112900
rect 197380 112880 197620 112900
rect 197880 112880 198120 112900
rect 198380 112880 198620 112900
rect 198880 112880 199120 112900
rect 199380 112880 199620 112900
rect 199880 112880 200120 112900
rect 200380 112880 200620 112900
rect 200880 112880 201120 112900
rect 201380 112880 201620 112900
rect 201880 112880 202120 112900
rect 202380 112880 202620 112900
rect 202880 112880 203120 112900
rect 203380 112880 203620 112900
rect 203880 112880 204120 112900
rect 204380 112880 204620 112900
rect 204880 112880 205120 112900
rect 205380 112880 205620 112900
rect 205880 112880 206120 112900
rect 206380 112880 206620 112900
rect 206880 112880 207120 112900
rect 207380 112880 207620 112900
rect 207880 112880 208120 112900
rect 208380 112880 208620 112900
rect 208880 112880 209120 112900
rect 209380 112880 209620 112900
rect 209880 112880 210120 112900
rect 210380 112880 210620 112900
rect 210880 112880 211120 112900
rect 211380 112880 211620 112900
rect 211880 112880 212120 112900
rect 212380 112880 212620 112900
rect 212880 112880 213120 112900
rect 213380 112880 213620 112900
rect 213880 112880 214120 112900
rect 214380 112880 214620 112900
rect 214880 112880 215120 112900
rect 215380 112880 215620 112900
rect 215880 112880 216120 112900
rect 216380 112880 216620 112900
rect 216880 112880 217120 112900
rect 217380 112880 217620 112900
rect 217880 112880 218120 112900
rect 218380 112880 218620 112900
rect 218880 112880 219120 112900
rect 219380 112880 219620 112900
rect 219880 112880 220120 112900
rect 220380 112880 220620 112900
rect 220880 112880 221120 112900
rect 221380 112880 221620 112900
rect 221880 112880 222120 112900
rect 222380 112880 222620 112900
rect 222880 112880 223120 112900
rect 223380 112880 223620 112900
rect 223880 112880 224120 112900
rect 224380 112880 224620 112900
rect 224880 112880 225120 112900
rect 225380 112880 225620 112900
rect 225880 112880 226120 112900
rect 226380 112880 226620 112900
rect 226880 112880 227120 112900
rect 227380 112880 227620 112900
rect 227880 112880 228120 112900
rect 228380 112880 228620 112900
rect 228880 112880 229120 112900
rect 229380 112880 229620 112900
rect 229880 112880 230120 112900
rect 230380 112880 230620 112900
rect 230880 112880 231120 112900
rect 231380 112880 231620 112900
rect 231880 112880 232000 112900
rect 178000 112620 178100 112880
rect 178400 112620 178600 112880
rect 178900 112620 179100 112880
rect 179400 112620 179600 112880
rect 179900 112620 180100 112880
rect 180400 112620 180600 112880
rect 180900 112620 181100 112880
rect 181400 112620 181600 112880
rect 181900 112620 182100 112880
rect 182400 112620 182600 112880
rect 182900 112620 183100 112880
rect 183400 112620 183600 112880
rect 183900 112620 184100 112880
rect 184400 112620 184600 112880
rect 184900 112620 185100 112880
rect 185400 112620 185600 112880
rect 185900 112620 186100 112880
rect 186400 112620 186600 112880
rect 186900 112620 187100 112880
rect 187400 112620 187600 112880
rect 187900 112620 188100 112880
rect 188400 112620 188600 112880
rect 188900 112620 189100 112880
rect 189400 112620 189600 112880
rect 189900 112620 190100 112880
rect 190400 112620 190600 112880
rect 190900 112620 191100 112880
rect 191400 112620 191600 112880
rect 191900 112620 192100 112880
rect 192400 112620 192600 112880
rect 192900 112620 193100 112880
rect 193400 112620 193600 112880
rect 193900 112620 194100 112880
rect 194400 112620 194600 112880
rect 194900 112620 195100 112880
rect 195400 112620 195600 112880
rect 195900 112620 196100 112880
rect 196400 112620 196600 112880
rect 196900 112620 197100 112880
rect 197400 112620 197600 112880
rect 197900 112620 198100 112880
rect 198400 112620 198600 112880
rect 198900 112620 199100 112880
rect 199400 112620 199600 112880
rect 199900 112620 200100 112880
rect 200400 112620 200600 112880
rect 200900 112620 201100 112880
rect 201400 112620 201600 112880
rect 201900 112620 202100 112880
rect 202400 112620 202600 112880
rect 202900 112620 203100 112880
rect 203400 112620 203600 112880
rect 203900 112620 204100 112880
rect 204400 112620 204600 112880
rect 204900 112620 205100 112880
rect 205400 112620 205600 112880
rect 205900 112620 206100 112880
rect 206400 112620 206600 112880
rect 206900 112620 207100 112880
rect 207400 112620 207600 112880
rect 207900 112620 208100 112880
rect 208400 112620 208600 112880
rect 208900 112620 209100 112880
rect 209400 112620 209600 112880
rect 209900 112620 210100 112880
rect 210400 112620 210600 112880
rect 210900 112620 211100 112880
rect 211400 112620 211600 112880
rect 211900 112620 212100 112880
rect 212400 112620 212600 112880
rect 212900 112620 213100 112880
rect 213400 112620 213600 112880
rect 213900 112620 214100 112880
rect 214400 112620 214600 112880
rect 214900 112620 215100 112880
rect 215400 112620 215600 112880
rect 215900 112620 216100 112880
rect 216400 112620 216600 112880
rect 216900 112620 217100 112880
rect 217400 112620 217600 112880
rect 217900 112620 218100 112880
rect 218400 112620 218600 112880
rect 218900 112620 219100 112880
rect 219400 112620 219600 112880
rect 219900 112620 220100 112880
rect 220400 112620 220600 112880
rect 220900 112620 221100 112880
rect 221400 112620 221600 112880
rect 221900 112620 222100 112880
rect 222400 112620 222600 112880
rect 222900 112620 223100 112880
rect 223400 112620 223600 112880
rect 223900 112620 224100 112880
rect 224400 112620 224600 112880
rect 224900 112620 225100 112880
rect 225400 112620 225600 112880
rect 225900 112620 226100 112880
rect 226400 112620 226600 112880
rect 226900 112620 227100 112880
rect 227400 112620 227600 112880
rect 227900 112620 228100 112880
rect 228400 112620 228600 112880
rect 228900 112620 229100 112880
rect 229400 112620 229600 112880
rect 229900 112620 230100 112880
rect 230400 112620 230600 112880
rect 230900 112620 231100 112880
rect 231400 112620 231600 112880
rect 231900 112620 232000 112880
rect 178000 112600 178120 112620
rect 178380 112600 178620 112620
rect 178880 112600 179120 112620
rect 179380 112600 179620 112620
rect 179880 112600 180120 112620
rect 180380 112600 180620 112620
rect 180880 112600 181120 112620
rect 181380 112600 181620 112620
rect 181880 112600 182120 112620
rect 182380 112600 182620 112620
rect 182880 112600 183120 112620
rect 183380 112600 183620 112620
rect 183880 112600 184120 112620
rect 184380 112600 184620 112620
rect 184880 112600 185120 112620
rect 185380 112600 185620 112620
rect 185880 112600 186120 112620
rect 186380 112600 186620 112620
rect 186880 112600 187120 112620
rect 187380 112600 187620 112620
rect 187880 112600 188120 112620
rect 188380 112600 188620 112620
rect 188880 112600 189120 112620
rect 189380 112600 189620 112620
rect 189880 112600 190120 112620
rect 190380 112600 190620 112620
rect 190880 112600 191120 112620
rect 191380 112600 191620 112620
rect 191880 112600 192120 112620
rect 192380 112600 192620 112620
rect 192880 112600 193120 112620
rect 193380 112600 193620 112620
rect 193880 112600 194120 112620
rect 194380 112600 194620 112620
rect 194880 112600 195120 112620
rect 195380 112600 195620 112620
rect 195880 112600 196120 112620
rect 196380 112600 196620 112620
rect 196880 112600 197120 112620
rect 197380 112600 197620 112620
rect 197880 112600 198120 112620
rect 198380 112600 198620 112620
rect 198880 112600 199120 112620
rect 199380 112600 199620 112620
rect 199880 112600 200120 112620
rect 200380 112600 200620 112620
rect 200880 112600 201120 112620
rect 201380 112600 201620 112620
rect 201880 112600 202120 112620
rect 202380 112600 202620 112620
rect 202880 112600 203120 112620
rect 203380 112600 203620 112620
rect 203880 112600 204120 112620
rect 204380 112600 204620 112620
rect 204880 112600 205120 112620
rect 205380 112600 205620 112620
rect 205880 112600 206120 112620
rect 206380 112600 206620 112620
rect 206880 112600 207120 112620
rect 207380 112600 207620 112620
rect 207880 112600 208120 112620
rect 208380 112600 208620 112620
rect 208880 112600 209120 112620
rect 209380 112600 209620 112620
rect 209880 112600 210120 112620
rect 210380 112600 210620 112620
rect 210880 112600 211120 112620
rect 211380 112600 211620 112620
rect 211880 112600 212120 112620
rect 212380 112600 212620 112620
rect 212880 112600 213120 112620
rect 213380 112600 213620 112620
rect 213880 112600 214120 112620
rect 214380 112600 214620 112620
rect 214880 112600 215120 112620
rect 215380 112600 215620 112620
rect 215880 112600 216120 112620
rect 216380 112600 216620 112620
rect 216880 112600 217120 112620
rect 217380 112600 217620 112620
rect 217880 112600 218120 112620
rect 218380 112600 218620 112620
rect 218880 112600 219120 112620
rect 219380 112600 219620 112620
rect 219880 112600 220120 112620
rect 220380 112600 220620 112620
rect 220880 112600 221120 112620
rect 221380 112600 221620 112620
rect 221880 112600 222120 112620
rect 222380 112600 222620 112620
rect 222880 112600 223120 112620
rect 223380 112600 223620 112620
rect 223880 112600 224120 112620
rect 224380 112600 224620 112620
rect 224880 112600 225120 112620
rect 225380 112600 225620 112620
rect 225880 112600 226120 112620
rect 226380 112600 226620 112620
rect 226880 112600 227120 112620
rect 227380 112600 227620 112620
rect 227880 112600 228120 112620
rect 228380 112600 228620 112620
rect 228880 112600 229120 112620
rect 229380 112600 229620 112620
rect 229880 112600 230120 112620
rect 230380 112600 230620 112620
rect 230880 112600 231120 112620
rect 231380 112600 231620 112620
rect 231880 112600 232000 112620
rect 178000 112400 232000 112600
rect 178000 112380 178120 112400
rect 178380 112380 178620 112400
rect 178880 112380 179120 112400
rect 179380 112380 179620 112400
rect 179880 112380 180120 112400
rect 180380 112380 180620 112400
rect 180880 112380 181120 112400
rect 181380 112380 181620 112400
rect 181880 112380 182120 112400
rect 182380 112380 182620 112400
rect 182880 112380 183120 112400
rect 183380 112380 183620 112400
rect 183880 112380 184120 112400
rect 184380 112380 184620 112400
rect 184880 112380 185120 112400
rect 185380 112380 185620 112400
rect 185880 112380 186120 112400
rect 186380 112380 186620 112400
rect 186880 112380 187120 112400
rect 187380 112380 187620 112400
rect 187880 112380 188120 112400
rect 188380 112380 188620 112400
rect 188880 112380 189120 112400
rect 189380 112380 189620 112400
rect 189880 112380 190120 112400
rect 190380 112380 190620 112400
rect 190880 112380 191120 112400
rect 191380 112380 191620 112400
rect 191880 112380 192120 112400
rect 192380 112380 192620 112400
rect 192880 112380 193120 112400
rect 193380 112380 193620 112400
rect 193880 112380 194120 112400
rect 194380 112380 194620 112400
rect 194880 112380 195120 112400
rect 195380 112380 195620 112400
rect 195880 112380 196120 112400
rect 196380 112380 196620 112400
rect 196880 112380 197120 112400
rect 197380 112380 197620 112400
rect 197880 112380 198120 112400
rect 198380 112380 198620 112400
rect 198880 112380 199120 112400
rect 199380 112380 199620 112400
rect 199880 112380 200120 112400
rect 200380 112380 200620 112400
rect 200880 112380 201120 112400
rect 201380 112380 201620 112400
rect 201880 112380 202120 112400
rect 202380 112380 202620 112400
rect 202880 112380 203120 112400
rect 203380 112380 203620 112400
rect 203880 112380 204120 112400
rect 204380 112380 204620 112400
rect 204880 112380 205120 112400
rect 205380 112380 205620 112400
rect 205880 112380 206120 112400
rect 206380 112380 206620 112400
rect 206880 112380 207120 112400
rect 207380 112380 207620 112400
rect 207880 112380 208120 112400
rect 208380 112380 208620 112400
rect 208880 112380 209120 112400
rect 209380 112380 209620 112400
rect 209880 112380 210120 112400
rect 210380 112380 210620 112400
rect 210880 112380 211120 112400
rect 211380 112380 211620 112400
rect 211880 112380 212120 112400
rect 212380 112380 212620 112400
rect 212880 112380 213120 112400
rect 213380 112380 213620 112400
rect 213880 112380 214120 112400
rect 214380 112380 214620 112400
rect 214880 112380 215120 112400
rect 215380 112380 215620 112400
rect 215880 112380 216120 112400
rect 216380 112380 216620 112400
rect 216880 112380 217120 112400
rect 217380 112380 217620 112400
rect 217880 112380 218120 112400
rect 218380 112380 218620 112400
rect 218880 112380 219120 112400
rect 219380 112380 219620 112400
rect 219880 112380 220120 112400
rect 220380 112380 220620 112400
rect 220880 112380 221120 112400
rect 221380 112380 221620 112400
rect 221880 112380 222120 112400
rect 222380 112380 222620 112400
rect 222880 112380 223120 112400
rect 223380 112380 223620 112400
rect 223880 112380 224120 112400
rect 224380 112380 224620 112400
rect 224880 112380 225120 112400
rect 225380 112380 225620 112400
rect 225880 112380 226120 112400
rect 226380 112380 226620 112400
rect 226880 112380 227120 112400
rect 227380 112380 227620 112400
rect 227880 112380 228120 112400
rect 228380 112380 228620 112400
rect 228880 112380 229120 112400
rect 229380 112380 229620 112400
rect 229880 112380 230120 112400
rect 230380 112380 230620 112400
rect 230880 112380 231120 112400
rect 231380 112380 231620 112400
rect 231880 112380 232000 112400
rect 178000 112120 178100 112380
rect 178400 112120 178600 112380
rect 178900 112120 179100 112380
rect 179400 112120 179600 112380
rect 179900 112120 180100 112380
rect 180400 112120 180600 112380
rect 180900 112120 181100 112380
rect 181400 112120 181600 112380
rect 181900 112120 182100 112380
rect 182400 112120 182600 112380
rect 182900 112120 183100 112380
rect 183400 112120 183600 112380
rect 183900 112120 184100 112380
rect 184400 112120 184600 112380
rect 184900 112120 185100 112380
rect 185400 112120 185600 112380
rect 185900 112120 186100 112380
rect 186400 112120 186600 112380
rect 186900 112120 187100 112380
rect 187400 112120 187600 112380
rect 187900 112120 188100 112380
rect 188400 112120 188600 112380
rect 188900 112120 189100 112380
rect 189400 112120 189600 112380
rect 189900 112120 190100 112380
rect 190400 112120 190600 112380
rect 190900 112120 191100 112380
rect 191400 112120 191600 112380
rect 191900 112120 192100 112380
rect 192400 112120 192600 112380
rect 192900 112120 193100 112380
rect 193400 112120 193600 112380
rect 193900 112120 194100 112380
rect 194400 112120 194600 112380
rect 194900 112120 195100 112380
rect 195400 112120 195600 112380
rect 195900 112120 196100 112380
rect 196400 112120 196600 112380
rect 196900 112120 197100 112380
rect 197400 112120 197600 112380
rect 197900 112120 198100 112380
rect 198400 112120 198600 112380
rect 198900 112120 199100 112380
rect 199400 112120 199600 112380
rect 199900 112120 200100 112380
rect 200400 112120 200600 112380
rect 200900 112120 201100 112380
rect 201400 112120 201600 112380
rect 201900 112120 202100 112380
rect 202400 112120 202600 112380
rect 202900 112120 203100 112380
rect 203400 112120 203600 112380
rect 203900 112120 204100 112380
rect 204400 112120 204600 112380
rect 204900 112120 205100 112380
rect 205400 112120 205600 112380
rect 205900 112120 206100 112380
rect 206400 112120 206600 112380
rect 206900 112120 207100 112380
rect 207400 112120 207600 112380
rect 207900 112120 208100 112380
rect 208400 112120 208600 112380
rect 208900 112120 209100 112380
rect 209400 112120 209600 112380
rect 209900 112120 210100 112380
rect 210400 112120 210600 112380
rect 210900 112120 211100 112380
rect 211400 112120 211600 112380
rect 211900 112120 212100 112380
rect 212400 112120 212600 112380
rect 212900 112120 213100 112380
rect 213400 112120 213600 112380
rect 213900 112120 214100 112380
rect 214400 112120 214600 112380
rect 214900 112120 215100 112380
rect 215400 112120 215600 112380
rect 215900 112120 216100 112380
rect 216400 112120 216600 112380
rect 216900 112120 217100 112380
rect 217400 112120 217600 112380
rect 217900 112120 218100 112380
rect 218400 112120 218600 112380
rect 218900 112120 219100 112380
rect 219400 112120 219600 112380
rect 219900 112120 220100 112380
rect 220400 112120 220600 112380
rect 220900 112120 221100 112380
rect 221400 112120 221600 112380
rect 221900 112120 222100 112380
rect 222400 112120 222600 112380
rect 222900 112120 223100 112380
rect 223400 112120 223600 112380
rect 223900 112120 224100 112380
rect 224400 112120 224600 112380
rect 224900 112120 225100 112380
rect 225400 112120 225600 112380
rect 225900 112120 226100 112380
rect 226400 112120 226600 112380
rect 226900 112120 227100 112380
rect 227400 112120 227600 112380
rect 227900 112120 228100 112380
rect 228400 112120 228600 112380
rect 228900 112120 229100 112380
rect 229400 112120 229600 112380
rect 229900 112120 230100 112380
rect 230400 112120 230600 112380
rect 230900 112120 231100 112380
rect 231400 112120 231600 112380
rect 231900 112120 232000 112380
rect 178000 112100 178120 112120
rect 178380 112100 178620 112120
rect 178880 112100 179120 112120
rect 179380 112100 179620 112120
rect 179880 112100 180120 112120
rect 180380 112100 180620 112120
rect 180880 112100 181120 112120
rect 181380 112100 181620 112120
rect 181880 112100 182120 112120
rect 182380 112100 182620 112120
rect 182880 112100 183120 112120
rect 183380 112100 183620 112120
rect 183880 112100 184120 112120
rect 184380 112100 184620 112120
rect 184880 112100 185120 112120
rect 185380 112100 185620 112120
rect 185880 112100 186120 112120
rect 186380 112100 186620 112120
rect 186880 112100 187120 112120
rect 187380 112100 187620 112120
rect 187880 112100 188120 112120
rect 188380 112100 188620 112120
rect 188880 112100 189120 112120
rect 189380 112100 189620 112120
rect 189880 112100 190120 112120
rect 190380 112100 190620 112120
rect 190880 112100 191120 112120
rect 191380 112100 191620 112120
rect 191880 112100 192120 112120
rect 192380 112100 192620 112120
rect 192880 112100 193120 112120
rect 193380 112100 193620 112120
rect 193880 112100 194120 112120
rect 194380 112100 194620 112120
rect 194880 112100 195120 112120
rect 195380 112100 195620 112120
rect 195880 112100 196120 112120
rect 196380 112100 196620 112120
rect 196880 112100 197120 112120
rect 197380 112100 197620 112120
rect 197880 112100 198120 112120
rect 198380 112100 198620 112120
rect 198880 112100 199120 112120
rect 199380 112100 199620 112120
rect 199880 112100 200120 112120
rect 200380 112100 200620 112120
rect 200880 112100 201120 112120
rect 201380 112100 201620 112120
rect 201880 112100 202120 112120
rect 202380 112100 202620 112120
rect 202880 112100 203120 112120
rect 203380 112100 203620 112120
rect 203880 112100 204120 112120
rect 204380 112100 204620 112120
rect 204880 112100 205120 112120
rect 205380 112100 205620 112120
rect 205880 112100 206120 112120
rect 206380 112100 206620 112120
rect 206880 112100 207120 112120
rect 207380 112100 207620 112120
rect 207880 112100 208120 112120
rect 208380 112100 208620 112120
rect 208880 112100 209120 112120
rect 209380 112100 209620 112120
rect 209880 112100 210120 112120
rect 210380 112100 210620 112120
rect 210880 112100 211120 112120
rect 211380 112100 211620 112120
rect 211880 112100 212120 112120
rect 212380 112100 212620 112120
rect 212880 112100 213120 112120
rect 213380 112100 213620 112120
rect 213880 112100 214120 112120
rect 214380 112100 214620 112120
rect 214880 112100 215120 112120
rect 215380 112100 215620 112120
rect 215880 112100 216120 112120
rect 216380 112100 216620 112120
rect 216880 112100 217120 112120
rect 217380 112100 217620 112120
rect 217880 112100 218120 112120
rect 218380 112100 218620 112120
rect 218880 112100 219120 112120
rect 219380 112100 219620 112120
rect 219880 112100 220120 112120
rect 220380 112100 220620 112120
rect 220880 112100 221120 112120
rect 221380 112100 221620 112120
rect 221880 112100 222120 112120
rect 222380 112100 222620 112120
rect 222880 112100 223120 112120
rect 223380 112100 223620 112120
rect 223880 112100 224120 112120
rect 224380 112100 224620 112120
rect 224880 112100 225120 112120
rect 225380 112100 225620 112120
rect 225880 112100 226120 112120
rect 226380 112100 226620 112120
rect 226880 112100 227120 112120
rect 227380 112100 227620 112120
rect 227880 112100 228120 112120
rect 228380 112100 228620 112120
rect 228880 112100 229120 112120
rect 229380 112100 229620 112120
rect 229880 112100 230120 112120
rect 230380 112100 230620 112120
rect 230880 112100 231120 112120
rect 231380 112100 231620 112120
rect 231880 112100 232000 112120
rect 178000 111900 232000 112100
rect 178000 111880 178120 111900
rect 178380 111880 178620 111900
rect 178880 111880 179120 111900
rect 179380 111880 179620 111900
rect 179880 111880 180120 111900
rect 180380 111880 180620 111900
rect 180880 111880 181120 111900
rect 181380 111880 181620 111900
rect 181880 111880 182120 111900
rect 182380 111880 182620 111900
rect 182880 111880 183120 111900
rect 183380 111880 183620 111900
rect 183880 111880 184120 111900
rect 184380 111880 184620 111900
rect 184880 111880 185120 111900
rect 185380 111880 185620 111900
rect 185880 111880 186120 111900
rect 186380 111880 186620 111900
rect 186880 111880 187120 111900
rect 187380 111880 187620 111900
rect 187880 111880 188120 111900
rect 188380 111880 188620 111900
rect 188880 111880 189120 111900
rect 189380 111880 189620 111900
rect 189880 111880 190120 111900
rect 190380 111880 190620 111900
rect 190880 111880 191120 111900
rect 191380 111880 191620 111900
rect 191880 111880 192120 111900
rect 192380 111880 192620 111900
rect 192880 111880 193120 111900
rect 193380 111880 193620 111900
rect 193880 111880 194120 111900
rect 194380 111880 194620 111900
rect 194880 111880 195120 111900
rect 195380 111880 195620 111900
rect 195880 111880 196120 111900
rect 196380 111880 196620 111900
rect 196880 111880 197120 111900
rect 197380 111880 197620 111900
rect 197880 111880 198120 111900
rect 198380 111880 198620 111900
rect 198880 111880 199120 111900
rect 199380 111880 199620 111900
rect 199880 111880 200120 111900
rect 200380 111880 200620 111900
rect 200880 111880 201120 111900
rect 201380 111880 201620 111900
rect 201880 111880 202120 111900
rect 202380 111880 202620 111900
rect 202880 111880 203120 111900
rect 203380 111880 203620 111900
rect 203880 111880 204120 111900
rect 204380 111880 204620 111900
rect 204880 111880 205120 111900
rect 205380 111880 205620 111900
rect 205880 111880 206120 111900
rect 206380 111880 206620 111900
rect 206880 111880 207120 111900
rect 207380 111880 207620 111900
rect 207880 111880 208120 111900
rect 208380 111880 208620 111900
rect 208880 111880 209120 111900
rect 209380 111880 209620 111900
rect 209880 111880 210120 111900
rect 210380 111880 210620 111900
rect 210880 111880 211120 111900
rect 211380 111880 211620 111900
rect 211880 111880 212120 111900
rect 212380 111880 212620 111900
rect 212880 111880 213120 111900
rect 213380 111880 213620 111900
rect 213880 111880 214120 111900
rect 214380 111880 214620 111900
rect 214880 111880 215120 111900
rect 215380 111880 215620 111900
rect 215880 111880 216120 111900
rect 216380 111880 216620 111900
rect 216880 111880 217120 111900
rect 217380 111880 217620 111900
rect 217880 111880 218120 111900
rect 218380 111880 218620 111900
rect 218880 111880 219120 111900
rect 219380 111880 219620 111900
rect 219880 111880 220120 111900
rect 220380 111880 220620 111900
rect 220880 111880 221120 111900
rect 221380 111880 221620 111900
rect 221880 111880 222120 111900
rect 222380 111880 222620 111900
rect 222880 111880 223120 111900
rect 223380 111880 223620 111900
rect 223880 111880 224120 111900
rect 224380 111880 224620 111900
rect 224880 111880 225120 111900
rect 225380 111880 225620 111900
rect 225880 111880 226120 111900
rect 226380 111880 226620 111900
rect 226880 111880 227120 111900
rect 227380 111880 227620 111900
rect 227880 111880 228120 111900
rect 228380 111880 228620 111900
rect 228880 111880 229120 111900
rect 229380 111880 229620 111900
rect 229880 111880 230120 111900
rect 230380 111880 230620 111900
rect 230880 111880 231120 111900
rect 231380 111880 231620 111900
rect 231880 111880 232000 111900
rect 178000 111620 178100 111880
rect 178400 111620 178600 111880
rect 178900 111620 179100 111880
rect 179400 111620 179600 111880
rect 179900 111620 180100 111880
rect 180400 111620 180600 111880
rect 180900 111620 181100 111880
rect 181400 111620 181600 111880
rect 181900 111620 182100 111880
rect 182400 111620 182600 111880
rect 182900 111620 183100 111880
rect 183400 111620 183600 111880
rect 183900 111620 184100 111880
rect 184400 111620 184600 111880
rect 184900 111620 185100 111880
rect 185400 111620 185600 111880
rect 185900 111620 186100 111880
rect 186400 111620 186600 111880
rect 186900 111620 187100 111880
rect 187400 111620 187600 111880
rect 187900 111620 188100 111880
rect 188400 111620 188600 111880
rect 188900 111620 189100 111880
rect 189400 111620 189600 111880
rect 189900 111620 190100 111880
rect 190400 111620 190600 111880
rect 190900 111620 191100 111880
rect 191400 111620 191600 111880
rect 191900 111620 192100 111880
rect 192400 111620 192600 111880
rect 192900 111620 193100 111880
rect 193400 111620 193600 111880
rect 193900 111620 194100 111880
rect 194400 111620 194600 111880
rect 194900 111620 195100 111880
rect 195400 111620 195600 111880
rect 195900 111620 196100 111880
rect 196400 111620 196600 111880
rect 196900 111620 197100 111880
rect 197400 111620 197600 111880
rect 197900 111620 198100 111880
rect 198400 111620 198600 111880
rect 198900 111620 199100 111880
rect 199400 111620 199600 111880
rect 199900 111620 200100 111880
rect 200400 111620 200600 111880
rect 200900 111620 201100 111880
rect 201400 111620 201600 111880
rect 201900 111620 202100 111880
rect 202400 111620 202600 111880
rect 202900 111620 203100 111880
rect 203400 111620 203600 111880
rect 203900 111620 204100 111880
rect 204400 111620 204600 111880
rect 204900 111620 205100 111880
rect 205400 111620 205600 111880
rect 205900 111620 206100 111880
rect 206400 111620 206600 111880
rect 206900 111620 207100 111880
rect 207400 111620 207600 111880
rect 207900 111620 208100 111880
rect 208400 111620 208600 111880
rect 208900 111620 209100 111880
rect 209400 111620 209600 111880
rect 209900 111620 210100 111880
rect 210400 111620 210600 111880
rect 210900 111620 211100 111880
rect 211400 111620 211600 111880
rect 211900 111620 212100 111880
rect 212400 111620 212600 111880
rect 212900 111620 213100 111880
rect 213400 111620 213600 111880
rect 213900 111620 214100 111880
rect 214400 111620 214600 111880
rect 214900 111620 215100 111880
rect 215400 111620 215600 111880
rect 215900 111620 216100 111880
rect 216400 111620 216600 111880
rect 216900 111620 217100 111880
rect 217400 111620 217600 111880
rect 217900 111620 218100 111880
rect 218400 111620 218600 111880
rect 218900 111620 219100 111880
rect 219400 111620 219600 111880
rect 219900 111620 220100 111880
rect 220400 111620 220600 111880
rect 220900 111620 221100 111880
rect 221400 111620 221600 111880
rect 221900 111620 222100 111880
rect 222400 111620 222600 111880
rect 222900 111620 223100 111880
rect 223400 111620 223600 111880
rect 223900 111620 224100 111880
rect 224400 111620 224600 111880
rect 224900 111620 225100 111880
rect 225400 111620 225600 111880
rect 225900 111620 226100 111880
rect 226400 111620 226600 111880
rect 226900 111620 227100 111880
rect 227400 111620 227600 111880
rect 227900 111620 228100 111880
rect 228400 111620 228600 111880
rect 228900 111620 229100 111880
rect 229400 111620 229600 111880
rect 229900 111620 230100 111880
rect 230400 111620 230600 111880
rect 230900 111620 231100 111880
rect 231400 111620 231600 111880
rect 231900 111620 232000 111880
rect 178000 111600 178120 111620
rect 178380 111600 178620 111620
rect 178880 111600 179120 111620
rect 179380 111600 179620 111620
rect 179880 111600 180120 111620
rect 180380 111600 180620 111620
rect 180880 111600 181120 111620
rect 181380 111600 181620 111620
rect 181880 111600 182120 111620
rect 182380 111600 182620 111620
rect 182880 111600 183120 111620
rect 183380 111600 183620 111620
rect 183880 111600 184120 111620
rect 184380 111600 184620 111620
rect 184880 111600 185120 111620
rect 185380 111600 185620 111620
rect 185880 111600 186120 111620
rect 186380 111600 186620 111620
rect 186880 111600 187120 111620
rect 187380 111600 187620 111620
rect 187880 111600 188120 111620
rect 188380 111600 188620 111620
rect 188880 111600 189120 111620
rect 189380 111600 189620 111620
rect 189880 111600 190120 111620
rect 190380 111600 190620 111620
rect 190880 111600 191120 111620
rect 191380 111600 191620 111620
rect 191880 111600 192120 111620
rect 192380 111600 192620 111620
rect 192880 111600 193120 111620
rect 193380 111600 193620 111620
rect 193880 111600 194120 111620
rect 194380 111600 194620 111620
rect 194880 111600 195120 111620
rect 195380 111600 195620 111620
rect 195880 111600 196120 111620
rect 196380 111600 196620 111620
rect 196880 111600 197120 111620
rect 197380 111600 197620 111620
rect 197880 111600 198120 111620
rect 198380 111600 198620 111620
rect 198880 111600 199120 111620
rect 199380 111600 199620 111620
rect 199880 111600 200120 111620
rect 200380 111600 200620 111620
rect 200880 111600 201120 111620
rect 201380 111600 201620 111620
rect 201880 111600 202120 111620
rect 202380 111600 202620 111620
rect 202880 111600 203120 111620
rect 203380 111600 203620 111620
rect 203880 111600 204120 111620
rect 204380 111600 204620 111620
rect 204880 111600 205120 111620
rect 205380 111600 205620 111620
rect 205880 111600 206120 111620
rect 206380 111600 206620 111620
rect 206880 111600 207120 111620
rect 207380 111600 207620 111620
rect 207880 111600 208120 111620
rect 208380 111600 208620 111620
rect 208880 111600 209120 111620
rect 209380 111600 209620 111620
rect 209880 111600 210120 111620
rect 210380 111600 210620 111620
rect 210880 111600 211120 111620
rect 211380 111600 211620 111620
rect 211880 111600 212120 111620
rect 212380 111600 212620 111620
rect 212880 111600 213120 111620
rect 213380 111600 213620 111620
rect 213880 111600 214120 111620
rect 214380 111600 214620 111620
rect 214880 111600 215120 111620
rect 215380 111600 215620 111620
rect 215880 111600 216120 111620
rect 216380 111600 216620 111620
rect 216880 111600 217120 111620
rect 217380 111600 217620 111620
rect 217880 111600 218120 111620
rect 218380 111600 218620 111620
rect 218880 111600 219120 111620
rect 219380 111600 219620 111620
rect 219880 111600 220120 111620
rect 220380 111600 220620 111620
rect 220880 111600 221120 111620
rect 221380 111600 221620 111620
rect 221880 111600 222120 111620
rect 222380 111600 222620 111620
rect 222880 111600 223120 111620
rect 223380 111600 223620 111620
rect 223880 111600 224120 111620
rect 224380 111600 224620 111620
rect 224880 111600 225120 111620
rect 225380 111600 225620 111620
rect 225880 111600 226120 111620
rect 226380 111600 226620 111620
rect 226880 111600 227120 111620
rect 227380 111600 227620 111620
rect 227880 111600 228120 111620
rect 228380 111600 228620 111620
rect 228880 111600 229120 111620
rect 229380 111600 229620 111620
rect 229880 111600 230120 111620
rect 230380 111600 230620 111620
rect 230880 111600 231120 111620
rect 231380 111600 231620 111620
rect 231880 111600 232000 111620
rect 178000 111400 232000 111600
rect 178000 111380 178120 111400
rect 178380 111380 178620 111400
rect 178880 111380 179120 111400
rect 179380 111380 179620 111400
rect 179880 111380 180120 111400
rect 180380 111380 180620 111400
rect 180880 111380 181120 111400
rect 181380 111380 181620 111400
rect 181880 111380 182120 111400
rect 182380 111380 182620 111400
rect 182880 111380 183120 111400
rect 183380 111380 183620 111400
rect 183880 111380 184120 111400
rect 184380 111380 184620 111400
rect 184880 111380 185120 111400
rect 185380 111380 185620 111400
rect 185880 111380 186120 111400
rect 186380 111380 186620 111400
rect 186880 111380 187120 111400
rect 187380 111380 187620 111400
rect 187880 111380 188120 111400
rect 188380 111380 188620 111400
rect 188880 111380 189120 111400
rect 189380 111380 189620 111400
rect 189880 111380 190120 111400
rect 190380 111380 190620 111400
rect 190880 111380 191120 111400
rect 191380 111380 191620 111400
rect 191880 111380 192120 111400
rect 192380 111380 192620 111400
rect 192880 111380 193120 111400
rect 193380 111380 193620 111400
rect 193880 111380 194120 111400
rect 194380 111380 194620 111400
rect 194880 111380 195120 111400
rect 195380 111380 195620 111400
rect 195880 111380 196120 111400
rect 196380 111380 196620 111400
rect 196880 111380 197120 111400
rect 197380 111380 197620 111400
rect 197880 111380 198120 111400
rect 198380 111380 198620 111400
rect 198880 111380 199120 111400
rect 199380 111380 199620 111400
rect 199880 111380 200120 111400
rect 200380 111380 200620 111400
rect 200880 111380 201120 111400
rect 201380 111380 201620 111400
rect 201880 111380 202120 111400
rect 202380 111380 202620 111400
rect 202880 111380 203120 111400
rect 203380 111380 203620 111400
rect 203880 111380 204120 111400
rect 204380 111380 204620 111400
rect 204880 111380 205120 111400
rect 205380 111380 205620 111400
rect 205880 111380 206120 111400
rect 206380 111380 206620 111400
rect 206880 111380 207120 111400
rect 207380 111380 207620 111400
rect 207880 111380 208120 111400
rect 208380 111380 208620 111400
rect 208880 111380 209120 111400
rect 209380 111380 209620 111400
rect 209880 111380 210120 111400
rect 210380 111380 210620 111400
rect 210880 111380 211120 111400
rect 211380 111380 211620 111400
rect 211880 111380 212120 111400
rect 212380 111380 212620 111400
rect 212880 111380 213120 111400
rect 213380 111380 213620 111400
rect 213880 111380 214120 111400
rect 214380 111380 214620 111400
rect 214880 111380 215120 111400
rect 215380 111380 215620 111400
rect 215880 111380 216120 111400
rect 216380 111380 216620 111400
rect 216880 111380 217120 111400
rect 217380 111380 217620 111400
rect 217880 111380 218120 111400
rect 218380 111380 218620 111400
rect 218880 111380 219120 111400
rect 219380 111380 219620 111400
rect 219880 111380 220120 111400
rect 220380 111380 220620 111400
rect 220880 111380 221120 111400
rect 221380 111380 221620 111400
rect 221880 111380 222120 111400
rect 222380 111380 222620 111400
rect 222880 111380 223120 111400
rect 223380 111380 223620 111400
rect 223880 111380 224120 111400
rect 224380 111380 224620 111400
rect 224880 111380 225120 111400
rect 225380 111380 225620 111400
rect 225880 111380 226120 111400
rect 226380 111380 226620 111400
rect 226880 111380 227120 111400
rect 227380 111380 227620 111400
rect 227880 111380 228120 111400
rect 228380 111380 228620 111400
rect 228880 111380 229120 111400
rect 229380 111380 229620 111400
rect 229880 111380 230120 111400
rect 230380 111380 230620 111400
rect 230880 111380 231120 111400
rect 231380 111380 231620 111400
rect 231880 111380 232000 111400
rect 178000 111120 178100 111380
rect 178400 111120 178600 111380
rect 178900 111120 179100 111380
rect 179400 111120 179600 111380
rect 179900 111120 180100 111380
rect 180400 111120 180600 111380
rect 180900 111120 181100 111380
rect 181400 111120 181600 111380
rect 181900 111120 182100 111380
rect 182400 111120 182600 111380
rect 182900 111120 183100 111380
rect 183400 111120 183600 111380
rect 183900 111120 184100 111380
rect 184400 111120 184600 111380
rect 184900 111120 185100 111380
rect 185400 111120 185600 111380
rect 185900 111120 186100 111380
rect 186400 111120 186600 111380
rect 186900 111120 187100 111380
rect 187400 111120 187600 111380
rect 187900 111120 188100 111380
rect 188400 111120 188600 111380
rect 188900 111120 189100 111380
rect 189400 111120 189600 111380
rect 189900 111120 190100 111380
rect 190400 111120 190600 111380
rect 190900 111120 191100 111380
rect 191400 111120 191600 111380
rect 191900 111120 192100 111380
rect 192400 111120 192600 111380
rect 192900 111120 193100 111380
rect 193400 111120 193600 111380
rect 193900 111120 194100 111380
rect 194400 111120 194600 111380
rect 194900 111120 195100 111380
rect 195400 111120 195600 111380
rect 195900 111120 196100 111380
rect 196400 111120 196600 111380
rect 196900 111120 197100 111380
rect 197400 111120 197600 111380
rect 197900 111120 198100 111380
rect 198400 111120 198600 111380
rect 198900 111120 199100 111380
rect 199400 111120 199600 111380
rect 199900 111120 200100 111380
rect 200400 111120 200600 111380
rect 200900 111120 201100 111380
rect 201400 111120 201600 111380
rect 201900 111120 202100 111380
rect 202400 111120 202600 111380
rect 202900 111120 203100 111380
rect 203400 111120 203600 111380
rect 203900 111120 204100 111380
rect 204400 111120 204600 111380
rect 204900 111120 205100 111380
rect 205400 111120 205600 111380
rect 205900 111120 206100 111380
rect 206400 111120 206600 111380
rect 206900 111120 207100 111380
rect 207400 111120 207600 111380
rect 207900 111120 208100 111380
rect 208400 111120 208600 111380
rect 208900 111120 209100 111380
rect 209400 111120 209600 111380
rect 209900 111120 210100 111380
rect 210400 111120 210600 111380
rect 210900 111120 211100 111380
rect 211400 111120 211600 111380
rect 211900 111120 212100 111380
rect 212400 111120 212600 111380
rect 212900 111120 213100 111380
rect 213400 111120 213600 111380
rect 213900 111120 214100 111380
rect 214400 111120 214600 111380
rect 214900 111120 215100 111380
rect 215400 111120 215600 111380
rect 215900 111120 216100 111380
rect 216400 111120 216600 111380
rect 216900 111120 217100 111380
rect 217400 111120 217600 111380
rect 217900 111120 218100 111380
rect 218400 111120 218600 111380
rect 218900 111120 219100 111380
rect 219400 111120 219600 111380
rect 219900 111120 220100 111380
rect 220400 111120 220600 111380
rect 220900 111120 221100 111380
rect 221400 111120 221600 111380
rect 221900 111120 222100 111380
rect 222400 111120 222600 111380
rect 222900 111120 223100 111380
rect 223400 111120 223600 111380
rect 223900 111120 224100 111380
rect 224400 111120 224600 111380
rect 224900 111120 225100 111380
rect 225400 111120 225600 111380
rect 225900 111120 226100 111380
rect 226400 111120 226600 111380
rect 226900 111120 227100 111380
rect 227400 111120 227600 111380
rect 227900 111120 228100 111380
rect 228400 111120 228600 111380
rect 228900 111120 229100 111380
rect 229400 111120 229600 111380
rect 229900 111120 230100 111380
rect 230400 111120 230600 111380
rect 230900 111120 231100 111380
rect 231400 111120 231600 111380
rect 231900 111120 232000 111380
rect 178000 111100 178120 111120
rect 178380 111100 178620 111120
rect 178880 111100 179120 111120
rect 179380 111100 179620 111120
rect 179880 111100 180120 111120
rect 180380 111100 180620 111120
rect 180880 111100 181120 111120
rect 181380 111100 181620 111120
rect 181880 111100 182120 111120
rect 182380 111100 182620 111120
rect 182880 111100 183120 111120
rect 183380 111100 183620 111120
rect 183880 111100 184120 111120
rect 184380 111100 184620 111120
rect 184880 111100 185120 111120
rect 185380 111100 185620 111120
rect 185880 111100 186120 111120
rect 186380 111100 186620 111120
rect 186880 111100 187120 111120
rect 187380 111100 187620 111120
rect 187880 111100 188120 111120
rect 188380 111100 188620 111120
rect 188880 111100 189120 111120
rect 189380 111100 189620 111120
rect 189880 111100 190120 111120
rect 190380 111100 190620 111120
rect 190880 111100 191120 111120
rect 191380 111100 191620 111120
rect 191880 111100 192120 111120
rect 192380 111100 192620 111120
rect 192880 111100 193120 111120
rect 193380 111100 193620 111120
rect 193880 111100 194120 111120
rect 194380 111100 194620 111120
rect 194880 111100 195120 111120
rect 195380 111100 195620 111120
rect 195880 111100 196120 111120
rect 196380 111100 196620 111120
rect 196880 111100 197120 111120
rect 197380 111100 197620 111120
rect 197880 111100 198120 111120
rect 198380 111100 198620 111120
rect 198880 111100 199120 111120
rect 199380 111100 199620 111120
rect 199880 111100 200120 111120
rect 200380 111100 200620 111120
rect 200880 111100 201120 111120
rect 201380 111100 201620 111120
rect 201880 111100 202120 111120
rect 202380 111100 202620 111120
rect 202880 111100 203120 111120
rect 203380 111100 203620 111120
rect 203880 111100 204120 111120
rect 204380 111100 204620 111120
rect 204880 111100 205120 111120
rect 205380 111100 205620 111120
rect 205880 111100 206120 111120
rect 206380 111100 206620 111120
rect 206880 111100 207120 111120
rect 207380 111100 207620 111120
rect 207880 111100 208120 111120
rect 208380 111100 208620 111120
rect 208880 111100 209120 111120
rect 209380 111100 209620 111120
rect 209880 111100 210120 111120
rect 210380 111100 210620 111120
rect 210880 111100 211120 111120
rect 211380 111100 211620 111120
rect 211880 111100 212120 111120
rect 212380 111100 212620 111120
rect 212880 111100 213120 111120
rect 213380 111100 213620 111120
rect 213880 111100 214120 111120
rect 214380 111100 214620 111120
rect 214880 111100 215120 111120
rect 215380 111100 215620 111120
rect 215880 111100 216120 111120
rect 216380 111100 216620 111120
rect 216880 111100 217120 111120
rect 217380 111100 217620 111120
rect 217880 111100 218120 111120
rect 218380 111100 218620 111120
rect 218880 111100 219120 111120
rect 219380 111100 219620 111120
rect 219880 111100 220120 111120
rect 220380 111100 220620 111120
rect 220880 111100 221120 111120
rect 221380 111100 221620 111120
rect 221880 111100 222120 111120
rect 222380 111100 222620 111120
rect 222880 111100 223120 111120
rect 223380 111100 223620 111120
rect 223880 111100 224120 111120
rect 224380 111100 224620 111120
rect 224880 111100 225120 111120
rect 225380 111100 225620 111120
rect 225880 111100 226120 111120
rect 226380 111100 226620 111120
rect 226880 111100 227120 111120
rect 227380 111100 227620 111120
rect 227880 111100 228120 111120
rect 228380 111100 228620 111120
rect 228880 111100 229120 111120
rect 229380 111100 229620 111120
rect 229880 111100 230120 111120
rect 230380 111100 230620 111120
rect 230880 111100 231120 111120
rect 231380 111100 231620 111120
rect 231880 111100 232000 111120
rect 178000 110900 232000 111100
rect 178000 110880 178120 110900
rect 178380 110880 178620 110900
rect 178880 110880 179120 110900
rect 179380 110880 179620 110900
rect 179880 110880 180120 110900
rect 180380 110880 180620 110900
rect 180880 110880 181120 110900
rect 181380 110880 181620 110900
rect 181880 110880 182120 110900
rect 182380 110880 182620 110900
rect 182880 110880 183120 110900
rect 183380 110880 183620 110900
rect 183880 110880 184120 110900
rect 184380 110880 184620 110900
rect 184880 110880 185120 110900
rect 185380 110880 185620 110900
rect 185880 110880 186120 110900
rect 186380 110880 186620 110900
rect 186880 110880 187120 110900
rect 187380 110880 187620 110900
rect 187880 110880 188120 110900
rect 188380 110880 188620 110900
rect 188880 110880 189120 110900
rect 189380 110880 189620 110900
rect 189880 110880 190120 110900
rect 190380 110880 190620 110900
rect 190880 110880 191120 110900
rect 191380 110880 191620 110900
rect 191880 110880 192120 110900
rect 192380 110880 192620 110900
rect 192880 110880 193120 110900
rect 193380 110880 193620 110900
rect 193880 110880 194120 110900
rect 194380 110880 194620 110900
rect 194880 110880 195120 110900
rect 195380 110880 195620 110900
rect 195880 110880 196120 110900
rect 196380 110880 196620 110900
rect 196880 110880 197120 110900
rect 197380 110880 197620 110900
rect 197880 110880 198120 110900
rect 198380 110880 198620 110900
rect 198880 110880 199120 110900
rect 199380 110880 199620 110900
rect 199880 110880 200120 110900
rect 200380 110880 200620 110900
rect 200880 110880 201120 110900
rect 201380 110880 201620 110900
rect 201880 110880 202120 110900
rect 202380 110880 202620 110900
rect 202880 110880 203120 110900
rect 203380 110880 203620 110900
rect 203880 110880 204120 110900
rect 204380 110880 204620 110900
rect 204880 110880 205120 110900
rect 205380 110880 205620 110900
rect 205880 110880 206120 110900
rect 206380 110880 206620 110900
rect 206880 110880 207120 110900
rect 207380 110880 207620 110900
rect 207880 110880 208120 110900
rect 208380 110880 208620 110900
rect 208880 110880 209120 110900
rect 209380 110880 209620 110900
rect 209880 110880 210120 110900
rect 210380 110880 210620 110900
rect 210880 110880 211120 110900
rect 211380 110880 211620 110900
rect 211880 110880 212120 110900
rect 212380 110880 212620 110900
rect 212880 110880 213120 110900
rect 213380 110880 213620 110900
rect 213880 110880 214120 110900
rect 214380 110880 214620 110900
rect 214880 110880 215120 110900
rect 215380 110880 215620 110900
rect 215880 110880 216120 110900
rect 216380 110880 216620 110900
rect 216880 110880 217120 110900
rect 217380 110880 217620 110900
rect 217880 110880 218120 110900
rect 218380 110880 218620 110900
rect 218880 110880 219120 110900
rect 219380 110880 219620 110900
rect 219880 110880 220120 110900
rect 220380 110880 220620 110900
rect 220880 110880 221120 110900
rect 221380 110880 221620 110900
rect 221880 110880 222120 110900
rect 222380 110880 222620 110900
rect 222880 110880 223120 110900
rect 223380 110880 223620 110900
rect 223880 110880 224120 110900
rect 224380 110880 224620 110900
rect 224880 110880 225120 110900
rect 225380 110880 225620 110900
rect 225880 110880 226120 110900
rect 226380 110880 226620 110900
rect 226880 110880 227120 110900
rect 227380 110880 227620 110900
rect 227880 110880 228120 110900
rect 228380 110880 228620 110900
rect 228880 110880 229120 110900
rect 229380 110880 229620 110900
rect 229880 110880 230120 110900
rect 230380 110880 230620 110900
rect 230880 110880 231120 110900
rect 231380 110880 231620 110900
rect 231880 110880 232000 110900
rect 178000 110620 178100 110880
rect 178400 110620 178600 110880
rect 178900 110620 179100 110880
rect 179400 110620 179600 110880
rect 179900 110620 180100 110880
rect 180400 110620 180600 110880
rect 180900 110620 181100 110880
rect 181400 110620 181600 110880
rect 181900 110620 182100 110880
rect 182400 110620 182600 110880
rect 182900 110620 183100 110880
rect 183400 110620 183600 110880
rect 183900 110620 184100 110880
rect 184400 110620 184600 110880
rect 184900 110620 185100 110880
rect 185400 110620 185600 110880
rect 185900 110620 186100 110880
rect 186400 110620 186600 110880
rect 186900 110620 187100 110880
rect 187400 110620 187600 110880
rect 187900 110620 188100 110880
rect 188400 110620 188600 110880
rect 188900 110620 189100 110880
rect 189400 110620 189600 110880
rect 189900 110620 190100 110880
rect 190400 110620 190600 110880
rect 190900 110620 191100 110880
rect 191400 110620 191600 110880
rect 191900 110620 192100 110880
rect 192400 110620 192600 110880
rect 192900 110620 193100 110880
rect 193400 110620 193600 110880
rect 193900 110620 194100 110880
rect 194400 110620 194600 110880
rect 194900 110620 195100 110880
rect 195400 110620 195600 110880
rect 195900 110620 196100 110880
rect 196400 110620 196600 110880
rect 196900 110620 197100 110880
rect 197400 110620 197600 110880
rect 197900 110620 198100 110880
rect 198400 110620 198600 110880
rect 198900 110620 199100 110880
rect 199400 110620 199600 110880
rect 199900 110620 200100 110880
rect 200400 110620 200600 110880
rect 200900 110620 201100 110880
rect 201400 110620 201600 110880
rect 201900 110620 202100 110880
rect 202400 110620 202600 110880
rect 202900 110620 203100 110880
rect 203400 110620 203600 110880
rect 203900 110620 204100 110880
rect 204400 110620 204600 110880
rect 204900 110620 205100 110880
rect 205400 110620 205600 110880
rect 205900 110620 206100 110880
rect 206400 110620 206600 110880
rect 206900 110620 207100 110880
rect 207400 110620 207600 110880
rect 207900 110620 208100 110880
rect 208400 110620 208600 110880
rect 208900 110620 209100 110880
rect 209400 110620 209600 110880
rect 209900 110620 210100 110880
rect 210400 110620 210600 110880
rect 210900 110620 211100 110880
rect 211400 110620 211600 110880
rect 211900 110620 212100 110880
rect 212400 110620 212600 110880
rect 212900 110620 213100 110880
rect 213400 110620 213600 110880
rect 213900 110620 214100 110880
rect 214400 110620 214600 110880
rect 214900 110620 215100 110880
rect 215400 110620 215600 110880
rect 215900 110620 216100 110880
rect 216400 110620 216600 110880
rect 216900 110620 217100 110880
rect 217400 110620 217600 110880
rect 217900 110620 218100 110880
rect 218400 110620 218600 110880
rect 218900 110620 219100 110880
rect 219400 110620 219600 110880
rect 219900 110620 220100 110880
rect 220400 110620 220600 110880
rect 220900 110620 221100 110880
rect 221400 110620 221600 110880
rect 221900 110620 222100 110880
rect 222400 110620 222600 110880
rect 222900 110620 223100 110880
rect 223400 110620 223600 110880
rect 223900 110620 224100 110880
rect 224400 110620 224600 110880
rect 224900 110620 225100 110880
rect 225400 110620 225600 110880
rect 225900 110620 226100 110880
rect 226400 110620 226600 110880
rect 226900 110620 227100 110880
rect 227400 110620 227600 110880
rect 227900 110620 228100 110880
rect 228400 110620 228600 110880
rect 228900 110620 229100 110880
rect 229400 110620 229600 110880
rect 229900 110620 230100 110880
rect 230400 110620 230600 110880
rect 230900 110620 231100 110880
rect 231400 110620 231600 110880
rect 231900 110620 232000 110880
rect 178000 110600 178120 110620
rect 178380 110600 178620 110620
rect 178880 110600 179120 110620
rect 179380 110600 179620 110620
rect 179880 110600 180120 110620
rect 180380 110600 180620 110620
rect 180880 110600 181120 110620
rect 181380 110600 181620 110620
rect 181880 110600 182120 110620
rect 182380 110600 182620 110620
rect 182880 110600 183120 110620
rect 183380 110600 183620 110620
rect 183880 110600 184120 110620
rect 184380 110600 184620 110620
rect 184880 110600 185120 110620
rect 185380 110600 185620 110620
rect 185880 110600 186120 110620
rect 186380 110600 186620 110620
rect 186880 110600 187120 110620
rect 187380 110600 187620 110620
rect 187880 110600 188120 110620
rect 188380 110600 188620 110620
rect 188880 110600 189120 110620
rect 189380 110600 189620 110620
rect 189880 110600 190120 110620
rect 190380 110600 190620 110620
rect 190880 110600 191120 110620
rect 191380 110600 191620 110620
rect 191880 110600 192120 110620
rect 192380 110600 192620 110620
rect 192880 110600 193120 110620
rect 193380 110600 193620 110620
rect 193880 110600 194120 110620
rect 194380 110600 194620 110620
rect 194880 110600 195120 110620
rect 195380 110600 195620 110620
rect 195880 110600 196120 110620
rect 196380 110600 196620 110620
rect 196880 110600 197120 110620
rect 197380 110600 197620 110620
rect 197880 110600 198120 110620
rect 198380 110600 198620 110620
rect 198880 110600 199120 110620
rect 199380 110600 199620 110620
rect 199880 110600 200120 110620
rect 200380 110600 200620 110620
rect 200880 110600 201120 110620
rect 201380 110600 201620 110620
rect 201880 110600 202120 110620
rect 202380 110600 202620 110620
rect 202880 110600 203120 110620
rect 203380 110600 203620 110620
rect 203880 110600 204120 110620
rect 204380 110600 204620 110620
rect 204880 110600 205120 110620
rect 205380 110600 205620 110620
rect 205880 110600 206120 110620
rect 206380 110600 206620 110620
rect 206880 110600 207120 110620
rect 207380 110600 207620 110620
rect 207880 110600 208120 110620
rect 208380 110600 208620 110620
rect 208880 110600 209120 110620
rect 209380 110600 209620 110620
rect 209880 110600 210120 110620
rect 210380 110600 210620 110620
rect 210880 110600 211120 110620
rect 211380 110600 211620 110620
rect 211880 110600 212120 110620
rect 212380 110600 212620 110620
rect 212880 110600 213120 110620
rect 213380 110600 213620 110620
rect 213880 110600 214120 110620
rect 214380 110600 214620 110620
rect 214880 110600 215120 110620
rect 215380 110600 215620 110620
rect 215880 110600 216120 110620
rect 216380 110600 216620 110620
rect 216880 110600 217120 110620
rect 217380 110600 217620 110620
rect 217880 110600 218120 110620
rect 218380 110600 218620 110620
rect 218880 110600 219120 110620
rect 219380 110600 219620 110620
rect 219880 110600 220120 110620
rect 220380 110600 220620 110620
rect 220880 110600 221120 110620
rect 221380 110600 221620 110620
rect 221880 110600 222120 110620
rect 222380 110600 222620 110620
rect 222880 110600 223120 110620
rect 223380 110600 223620 110620
rect 223880 110600 224120 110620
rect 224380 110600 224620 110620
rect 224880 110600 225120 110620
rect 225380 110600 225620 110620
rect 225880 110600 226120 110620
rect 226380 110600 226620 110620
rect 226880 110600 227120 110620
rect 227380 110600 227620 110620
rect 227880 110600 228120 110620
rect 228380 110600 228620 110620
rect 228880 110600 229120 110620
rect 229380 110600 229620 110620
rect 229880 110600 230120 110620
rect 230380 110600 230620 110620
rect 230880 110600 231120 110620
rect 231380 110600 231620 110620
rect 231880 110600 232000 110620
rect 178000 110400 232000 110600
rect 178000 110380 178120 110400
rect 178380 110380 178620 110400
rect 178880 110380 179120 110400
rect 179380 110380 179620 110400
rect 179880 110380 180120 110400
rect 180380 110380 180620 110400
rect 180880 110380 181120 110400
rect 181380 110380 181620 110400
rect 181880 110380 182120 110400
rect 182380 110380 182620 110400
rect 182880 110380 183120 110400
rect 183380 110380 183620 110400
rect 183880 110380 184120 110400
rect 184380 110380 184620 110400
rect 184880 110380 185120 110400
rect 185380 110380 185620 110400
rect 185880 110380 186120 110400
rect 186380 110380 186620 110400
rect 186880 110380 187120 110400
rect 187380 110380 187620 110400
rect 187880 110380 188120 110400
rect 188380 110380 188620 110400
rect 188880 110380 189120 110400
rect 189380 110380 189620 110400
rect 189880 110380 190120 110400
rect 190380 110380 190620 110400
rect 190880 110380 191120 110400
rect 191380 110380 191620 110400
rect 191880 110380 192120 110400
rect 192380 110380 192620 110400
rect 192880 110380 193120 110400
rect 193380 110380 193620 110400
rect 193880 110380 194120 110400
rect 194380 110380 194620 110400
rect 194880 110380 195120 110400
rect 195380 110380 195620 110400
rect 195880 110380 196120 110400
rect 196380 110380 196620 110400
rect 196880 110380 197120 110400
rect 197380 110380 197620 110400
rect 197880 110380 198120 110400
rect 198380 110380 198620 110400
rect 198880 110380 199120 110400
rect 199380 110380 199620 110400
rect 199880 110380 200120 110400
rect 200380 110380 200620 110400
rect 200880 110380 201120 110400
rect 201380 110380 201620 110400
rect 201880 110380 202120 110400
rect 202380 110380 202620 110400
rect 202880 110380 203120 110400
rect 203380 110380 203620 110400
rect 203880 110380 204120 110400
rect 204380 110380 204620 110400
rect 204880 110380 205120 110400
rect 205380 110380 205620 110400
rect 205880 110380 206120 110400
rect 206380 110380 206620 110400
rect 206880 110380 207120 110400
rect 207380 110380 207620 110400
rect 207880 110380 208120 110400
rect 208380 110380 208620 110400
rect 208880 110380 209120 110400
rect 209380 110380 209620 110400
rect 209880 110380 210120 110400
rect 210380 110380 210620 110400
rect 210880 110380 211120 110400
rect 211380 110380 211620 110400
rect 211880 110380 212120 110400
rect 212380 110380 212620 110400
rect 212880 110380 213120 110400
rect 213380 110380 213620 110400
rect 213880 110380 214120 110400
rect 214380 110380 214620 110400
rect 214880 110380 215120 110400
rect 215380 110380 215620 110400
rect 215880 110380 216120 110400
rect 216380 110380 216620 110400
rect 216880 110380 217120 110400
rect 217380 110380 217620 110400
rect 217880 110380 218120 110400
rect 218380 110380 218620 110400
rect 218880 110380 219120 110400
rect 219380 110380 219620 110400
rect 219880 110380 220120 110400
rect 220380 110380 220620 110400
rect 220880 110380 221120 110400
rect 221380 110380 221620 110400
rect 221880 110380 222120 110400
rect 222380 110380 222620 110400
rect 222880 110380 223120 110400
rect 223380 110380 223620 110400
rect 223880 110380 224120 110400
rect 224380 110380 224620 110400
rect 224880 110380 225120 110400
rect 225380 110380 225620 110400
rect 225880 110380 226120 110400
rect 226380 110380 226620 110400
rect 226880 110380 227120 110400
rect 227380 110380 227620 110400
rect 227880 110380 228120 110400
rect 228380 110380 228620 110400
rect 228880 110380 229120 110400
rect 229380 110380 229620 110400
rect 229880 110380 230120 110400
rect 230380 110380 230620 110400
rect 230880 110380 231120 110400
rect 231380 110380 231620 110400
rect 231880 110380 232000 110400
rect 178000 110120 178100 110380
rect 178400 110120 178600 110380
rect 178900 110120 179100 110380
rect 179400 110120 179600 110380
rect 179900 110120 180100 110380
rect 180400 110120 180600 110380
rect 180900 110120 181100 110380
rect 181400 110120 181600 110380
rect 181900 110120 182100 110380
rect 182400 110120 182600 110380
rect 182900 110120 183100 110380
rect 183400 110120 183600 110380
rect 183900 110120 184100 110380
rect 184400 110120 184600 110380
rect 184900 110120 185100 110380
rect 185400 110120 185600 110380
rect 185900 110120 186100 110380
rect 186400 110120 186600 110380
rect 186900 110120 187100 110380
rect 187400 110120 187600 110380
rect 187900 110120 188100 110380
rect 188400 110120 188600 110380
rect 188900 110120 189100 110380
rect 189400 110120 189600 110380
rect 189900 110120 190100 110380
rect 190400 110120 190600 110380
rect 190900 110120 191100 110380
rect 191400 110120 191600 110380
rect 191900 110120 192100 110380
rect 192400 110120 192600 110380
rect 192900 110120 193100 110380
rect 193400 110120 193600 110380
rect 193900 110120 194100 110380
rect 194400 110120 194600 110380
rect 194900 110120 195100 110380
rect 195400 110120 195600 110380
rect 195900 110120 196100 110380
rect 196400 110120 196600 110380
rect 196900 110120 197100 110380
rect 197400 110120 197600 110380
rect 197900 110120 198100 110380
rect 198400 110120 198600 110380
rect 198900 110120 199100 110380
rect 199400 110120 199600 110380
rect 199900 110120 200100 110380
rect 200400 110120 200600 110380
rect 200900 110120 201100 110380
rect 201400 110120 201600 110380
rect 201900 110120 202100 110380
rect 202400 110120 202600 110380
rect 202900 110120 203100 110380
rect 203400 110120 203600 110380
rect 203900 110120 204100 110380
rect 204400 110120 204600 110380
rect 204900 110120 205100 110380
rect 205400 110120 205600 110380
rect 205900 110120 206100 110380
rect 206400 110120 206600 110380
rect 206900 110120 207100 110380
rect 207400 110120 207600 110380
rect 207900 110120 208100 110380
rect 208400 110120 208600 110380
rect 208900 110120 209100 110380
rect 209400 110120 209600 110380
rect 209900 110120 210100 110380
rect 210400 110120 210600 110380
rect 210900 110120 211100 110380
rect 211400 110120 211600 110380
rect 211900 110120 212100 110380
rect 212400 110120 212600 110380
rect 212900 110120 213100 110380
rect 213400 110120 213600 110380
rect 213900 110120 214100 110380
rect 214400 110120 214600 110380
rect 214900 110120 215100 110380
rect 215400 110120 215600 110380
rect 215900 110120 216100 110380
rect 216400 110120 216600 110380
rect 216900 110120 217100 110380
rect 217400 110120 217600 110380
rect 217900 110120 218100 110380
rect 218400 110120 218600 110380
rect 218900 110120 219100 110380
rect 219400 110120 219600 110380
rect 219900 110120 220100 110380
rect 220400 110120 220600 110380
rect 220900 110120 221100 110380
rect 221400 110120 221600 110380
rect 221900 110120 222100 110380
rect 222400 110120 222600 110380
rect 222900 110120 223100 110380
rect 223400 110120 223600 110380
rect 223900 110120 224100 110380
rect 224400 110120 224600 110380
rect 224900 110120 225100 110380
rect 225400 110120 225600 110380
rect 225900 110120 226100 110380
rect 226400 110120 226600 110380
rect 226900 110120 227100 110380
rect 227400 110120 227600 110380
rect 227900 110120 228100 110380
rect 228400 110120 228600 110380
rect 228900 110120 229100 110380
rect 229400 110120 229600 110380
rect 229900 110120 230100 110380
rect 230400 110120 230600 110380
rect 230900 110120 231100 110380
rect 231400 110120 231600 110380
rect 231900 110120 232000 110380
rect 178000 110100 178120 110120
rect 178380 110100 178620 110120
rect 178880 110100 179120 110120
rect 179380 110100 179620 110120
rect 179880 110100 180120 110120
rect 180380 110100 180620 110120
rect 180880 110100 181120 110120
rect 181380 110100 181620 110120
rect 181880 110100 182120 110120
rect 182380 110100 182620 110120
rect 182880 110100 183120 110120
rect 183380 110100 183620 110120
rect 183880 110100 184120 110120
rect 184380 110100 184620 110120
rect 184880 110100 185120 110120
rect 185380 110100 185620 110120
rect 185880 110100 186120 110120
rect 186380 110100 186620 110120
rect 186880 110100 187120 110120
rect 187380 110100 187620 110120
rect 187880 110100 188120 110120
rect 188380 110100 188620 110120
rect 188880 110100 189120 110120
rect 189380 110100 189620 110120
rect 189880 110100 190120 110120
rect 190380 110100 190620 110120
rect 190880 110100 191120 110120
rect 191380 110100 191620 110120
rect 191880 110100 192120 110120
rect 192380 110100 192620 110120
rect 192880 110100 193120 110120
rect 193380 110100 193620 110120
rect 193880 110100 194120 110120
rect 194380 110100 194620 110120
rect 194880 110100 195120 110120
rect 195380 110100 195620 110120
rect 195880 110100 196120 110120
rect 196380 110100 196620 110120
rect 196880 110100 197120 110120
rect 197380 110100 197620 110120
rect 197880 110100 198120 110120
rect 198380 110100 198620 110120
rect 198880 110100 199120 110120
rect 199380 110100 199620 110120
rect 199880 110100 200120 110120
rect 200380 110100 200620 110120
rect 200880 110100 201120 110120
rect 201380 110100 201620 110120
rect 201880 110100 202120 110120
rect 202380 110100 202620 110120
rect 202880 110100 203120 110120
rect 203380 110100 203620 110120
rect 203880 110100 204120 110120
rect 204380 110100 204620 110120
rect 204880 110100 205120 110120
rect 205380 110100 205620 110120
rect 205880 110100 206120 110120
rect 206380 110100 206620 110120
rect 206880 110100 207120 110120
rect 207380 110100 207620 110120
rect 207880 110100 208120 110120
rect 208380 110100 208620 110120
rect 208880 110100 209120 110120
rect 209380 110100 209620 110120
rect 209880 110100 210120 110120
rect 210380 110100 210620 110120
rect 210880 110100 211120 110120
rect 211380 110100 211620 110120
rect 211880 110100 212120 110120
rect 212380 110100 212620 110120
rect 212880 110100 213120 110120
rect 213380 110100 213620 110120
rect 213880 110100 214120 110120
rect 214380 110100 214620 110120
rect 214880 110100 215120 110120
rect 215380 110100 215620 110120
rect 215880 110100 216120 110120
rect 216380 110100 216620 110120
rect 216880 110100 217120 110120
rect 217380 110100 217620 110120
rect 217880 110100 218120 110120
rect 218380 110100 218620 110120
rect 218880 110100 219120 110120
rect 219380 110100 219620 110120
rect 219880 110100 220120 110120
rect 220380 110100 220620 110120
rect 220880 110100 221120 110120
rect 221380 110100 221620 110120
rect 221880 110100 222120 110120
rect 222380 110100 222620 110120
rect 222880 110100 223120 110120
rect 223380 110100 223620 110120
rect 223880 110100 224120 110120
rect 224380 110100 224620 110120
rect 224880 110100 225120 110120
rect 225380 110100 225620 110120
rect 225880 110100 226120 110120
rect 226380 110100 226620 110120
rect 226880 110100 227120 110120
rect 227380 110100 227620 110120
rect 227880 110100 228120 110120
rect 228380 110100 228620 110120
rect 228880 110100 229120 110120
rect 229380 110100 229620 110120
rect 229880 110100 230120 110120
rect 230380 110100 230620 110120
rect 230880 110100 231120 110120
rect 231380 110100 231620 110120
rect 231880 110100 232000 110120
rect 178000 109900 232000 110100
rect 178000 109880 178120 109900
rect 178380 109880 178620 109900
rect 178880 109880 179120 109900
rect 179380 109880 179620 109900
rect 179880 109880 180120 109900
rect 180380 109880 180620 109900
rect 180880 109880 181120 109900
rect 181380 109880 181620 109900
rect 181880 109880 182120 109900
rect 182380 109880 182620 109900
rect 182880 109880 183120 109900
rect 183380 109880 183620 109900
rect 183880 109880 184120 109900
rect 184380 109880 184620 109900
rect 184880 109880 185120 109900
rect 185380 109880 185620 109900
rect 185880 109880 186120 109900
rect 186380 109880 186620 109900
rect 186880 109880 187120 109900
rect 187380 109880 187620 109900
rect 187880 109880 188120 109900
rect 188380 109880 188620 109900
rect 188880 109880 189120 109900
rect 189380 109880 189620 109900
rect 189880 109880 190120 109900
rect 190380 109880 190620 109900
rect 190880 109880 191120 109900
rect 191380 109880 191620 109900
rect 191880 109880 192120 109900
rect 192380 109880 192620 109900
rect 192880 109880 193120 109900
rect 193380 109880 193620 109900
rect 193880 109880 194120 109900
rect 194380 109880 194620 109900
rect 194880 109880 195120 109900
rect 195380 109880 195620 109900
rect 195880 109880 196120 109900
rect 196380 109880 196620 109900
rect 196880 109880 197120 109900
rect 197380 109880 197620 109900
rect 197880 109880 198120 109900
rect 198380 109880 198620 109900
rect 198880 109880 199120 109900
rect 199380 109880 199620 109900
rect 199880 109880 200120 109900
rect 200380 109880 200620 109900
rect 200880 109880 201120 109900
rect 201380 109880 201620 109900
rect 201880 109880 202120 109900
rect 202380 109880 202620 109900
rect 202880 109880 203120 109900
rect 203380 109880 203620 109900
rect 203880 109880 204120 109900
rect 204380 109880 204620 109900
rect 204880 109880 205120 109900
rect 205380 109880 205620 109900
rect 205880 109880 206120 109900
rect 206380 109880 206620 109900
rect 206880 109880 207120 109900
rect 207380 109880 207620 109900
rect 207880 109880 208120 109900
rect 208380 109880 208620 109900
rect 208880 109880 209120 109900
rect 209380 109880 209620 109900
rect 209880 109880 210120 109900
rect 210380 109880 210620 109900
rect 210880 109880 211120 109900
rect 211380 109880 211620 109900
rect 211880 109880 212120 109900
rect 212380 109880 212620 109900
rect 212880 109880 213120 109900
rect 213380 109880 213620 109900
rect 213880 109880 214120 109900
rect 214380 109880 214620 109900
rect 214880 109880 215120 109900
rect 215380 109880 215620 109900
rect 215880 109880 216120 109900
rect 216380 109880 216620 109900
rect 216880 109880 217120 109900
rect 217380 109880 217620 109900
rect 217880 109880 218120 109900
rect 218380 109880 218620 109900
rect 218880 109880 219120 109900
rect 219380 109880 219620 109900
rect 219880 109880 220120 109900
rect 220380 109880 220620 109900
rect 220880 109880 221120 109900
rect 221380 109880 221620 109900
rect 221880 109880 222120 109900
rect 222380 109880 222620 109900
rect 222880 109880 223120 109900
rect 223380 109880 223620 109900
rect 223880 109880 224120 109900
rect 224380 109880 224620 109900
rect 224880 109880 225120 109900
rect 225380 109880 225620 109900
rect 225880 109880 226120 109900
rect 226380 109880 226620 109900
rect 226880 109880 227120 109900
rect 227380 109880 227620 109900
rect 227880 109880 228120 109900
rect 228380 109880 228620 109900
rect 228880 109880 229120 109900
rect 229380 109880 229620 109900
rect 229880 109880 230120 109900
rect 230380 109880 230620 109900
rect 230880 109880 231120 109900
rect 231380 109880 231620 109900
rect 231880 109880 232000 109900
rect 178000 109620 178100 109880
rect 178400 109620 178600 109880
rect 178900 109620 179100 109880
rect 179400 109620 179600 109880
rect 179900 109620 180100 109880
rect 180400 109620 180600 109880
rect 180900 109620 181100 109880
rect 181400 109620 181600 109880
rect 181900 109620 182100 109880
rect 182400 109620 182600 109880
rect 182900 109620 183100 109880
rect 183400 109620 183600 109880
rect 183900 109620 184100 109880
rect 184400 109620 184600 109880
rect 184900 109620 185100 109880
rect 185400 109620 185600 109880
rect 185900 109620 186100 109880
rect 186400 109620 186600 109880
rect 186900 109620 187100 109880
rect 187400 109620 187600 109880
rect 187900 109620 188100 109880
rect 188400 109620 188600 109880
rect 188900 109620 189100 109880
rect 189400 109620 189600 109880
rect 189900 109620 190100 109880
rect 190400 109620 190600 109880
rect 190900 109620 191100 109880
rect 191400 109620 191600 109880
rect 191900 109620 192100 109880
rect 192400 109620 192600 109880
rect 192900 109620 193100 109880
rect 193400 109620 193600 109880
rect 193900 109620 194100 109880
rect 194400 109620 194600 109880
rect 194900 109620 195100 109880
rect 195400 109620 195600 109880
rect 195900 109620 196100 109880
rect 196400 109620 196600 109880
rect 196900 109620 197100 109880
rect 197400 109620 197600 109880
rect 197900 109620 198100 109880
rect 198400 109620 198600 109880
rect 198900 109620 199100 109880
rect 199400 109620 199600 109880
rect 199900 109620 200100 109880
rect 200400 109620 200600 109880
rect 200900 109620 201100 109880
rect 201400 109620 201600 109880
rect 201900 109620 202100 109880
rect 202400 109620 202600 109880
rect 202900 109620 203100 109880
rect 203400 109620 203600 109880
rect 203900 109620 204100 109880
rect 204400 109620 204600 109880
rect 204900 109620 205100 109880
rect 205400 109620 205600 109880
rect 205900 109620 206100 109880
rect 206400 109620 206600 109880
rect 206900 109620 207100 109880
rect 207400 109620 207600 109880
rect 207900 109620 208100 109880
rect 208400 109620 208600 109880
rect 208900 109620 209100 109880
rect 209400 109620 209600 109880
rect 209900 109620 210100 109880
rect 210400 109620 210600 109880
rect 210900 109620 211100 109880
rect 211400 109620 211600 109880
rect 211900 109620 212100 109880
rect 212400 109620 212600 109880
rect 212900 109620 213100 109880
rect 213400 109620 213600 109880
rect 213900 109620 214100 109880
rect 214400 109620 214600 109880
rect 214900 109620 215100 109880
rect 215400 109620 215600 109880
rect 215900 109620 216100 109880
rect 216400 109620 216600 109880
rect 216900 109620 217100 109880
rect 217400 109620 217600 109880
rect 217900 109620 218100 109880
rect 218400 109620 218600 109880
rect 218900 109620 219100 109880
rect 219400 109620 219600 109880
rect 219900 109620 220100 109880
rect 220400 109620 220600 109880
rect 220900 109620 221100 109880
rect 221400 109620 221600 109880
rect 221900 109620 222100 109880
rect 222400 109620 222600 109880
rect 222900 109620 223100 109880
rect 223400 109620 223600 109880
rect 223900 109620 224100 109880
rect 224400 109620 224600 109880
rect 224900 109620 225100 109880
rect 225400 109620 225600 109880
rect 225900 109620 226100 109880
rect 226400 109620 226600 109880
rect 226900 109620 227100 109880
rect 227400 109620 227600 109880
rect 227900 109620 228100 109880
rect 228400 109620 228600 109880
rect 228900 109620 229100 109880
rect 229400 109620 229600 109880
rect 229900 109620 230100 109880
rect 230400 109620 230600 109880
rect 230900 109620 231100 109880
rect 231400 109620 231600 109880
rect 231900 109620 232000 109880
rect 178000 109600 178120 109620
rect 178380 109600 178620 109620
rect 178880 109600 179120 109620
rect 179380 109600 179620 109620
rect 179880 109600 180120 109620
rect 180380 109600 180620 109620
rect 180880 109600 181120 109620
rect 181380 109600 181620 109620
rect 181880 109600 182120 109620
rect 182380 109600 182620 109620
rect 182880 109600 183120 109620
rect 183380 109600 183620 109620
rect 183880 109600 184120 109620
rect 184380 109600 184620 109620
rect 184880 109600 185120 109620
rect 185380 109600 185620 109620
rect 185880 109600 186120 109620
rect 186380 109600 186620 109620
rect 186880 109600 187120 109620
rect 187380 109600 187620 109620
rect 187880 109600 188120 109620
rect 188380 109600 188620 109620
rect 188880 109600 189120 109620
rect 189380 109600 189620 109620
rect 189880 109600 190120 109620
rect 190380 109600 190620 109620
rect 190880 109600 191120 109620
rect 191380 109600 191620 109620
rect 191880 109600 192120 109620
rect 192380 109600 192620 109620
rect 192880 109600 193120 109620
rect 193380 109600 193620 109620
rect 193880 109600 194120 109620
rect 194380 109600 194620 109620
rect 194880 109600 195120 109620
rect 195380 109600 195620 109620
rect 195880 109600 196120 109620
rect 196380 109600 196620 109620
rect 196880 109600 197120 109620
rect 197380 109600 197620 109620
rect 197880 109600 198120 109620
rect 198380 109600 198620 109620
rect 198880 109600 199120 109620
rect 199380 109600 199620 109620
rect 199880 109600 200120 109620
rect 200380 109600 200620 109620
rect 200880 109600 201120 109620
rect 201380 109600 201620 109620
rect 201880 109600 202120 109620
rect 202380 109600 202620 109620
rect 202880 109600 203120 109620
rect 203380 109600 203620 109620
rect 203880 109600 204120 109620
rect 204380 109600 204620 109620
rect 204880 109600 205120 109620
rect 205380 109600 205620 109620
rect 205880 109600 206120 109620
rect 206380 109600 206620 109620
rect 206880 109600 207120 109620
rect 207380 109600 207620 109620
rect 207880 109600 208120 109620
rect 208380 109600 208620 109620
rect 208880 109600 209120 109620
rect 209380 109600 209620 109620
rect 209880 109600 210120 109620
rect 210380 109600 210620 109620
rect 210880 109600 211120 109620
rect 211380 109600 211620 109620
rect 211880 109600 212120 109620
rect 212380 109600 212620 109620
rect 212880 109600 213120 109620
rect 213380 109600 213620 109620
rect 213880 109600 214120 109620
rect 214380 109600 214620 109620
rect 214880 109600 215120 109620
rect 215380 109600 215620 109620
rect 215880 109600 216120 109620
rect 216380 109600 216620 109620
rect 216880 109600 217120 109620
rect 217380 109600 217620 109620
rect 217880 109600 218120 109620
rect 218380 109600 218620 109620
rect 218880 109600 219120 109620
rect 219380 109600 219620 109620
rect 219880 109600 220120 109620
rect 220380 109600 220620 109620
rect 220880 109600 221120 109620
rect 221380 109600 221620 109620
rect 221880 109600 222120 109620
rect 222380 109600 222620 109620
rect 222880 109600 223120 109620
rect 223380 109600 223620 109620
rect 223880 109600 224120 109620
rect 224380 109600 224620 109620
rect 224880 109600 225120 109620
rect 225380 109600 225620 109620
rect 225880 109600 226120 109620
rect 226380 109600 226620 109620
rect 226880 109600 227120 109620
rect 227380 109600 227620 109620
rect 227880 109600 228120 109620
rect 228380 109600 228620 109620
rect 228880 109600 229120 109620
rect 229380 109600 229620 109620
rect 229880 109600 230120 109620
rect 230380 109600 230620 109620
rect 230880 109600 231120 109620
rect 231380 109600 231620 109620
rect 231880 109600 232000 109620
rect 178000 109400 232000 109600
rect 178000 109380 178120 109400
rect 178380 109380 178620 109400
rect 178880 109380 179120 109400
rect 179380 109380 179620 109400
rect 179880 109380 180120 109400
rect 180380 109380 180620 109400
rect 180880 109380 181120 109400
rect 181380 109380 181620 109400
rect 181880 109380 182120 109400
rect 182380 109380 182620 109400
rect 182880 109380 183120 109400
rect 183380 109380 183620 109400
rect 183880 109380 184120 109400
rect 184380 109380 184620 109400
rect 184880 109380 185120 109400
rect 185380 109380 185620 109400
rect 185880 109380 186120 109400
rect 186380 109380 186620 109400
rect 186880 109380 187120 109400
rect 187380 109380 187620 109400
rect 187880 109380 188120 109400
rect 188380 109380 188620 109400
rect 188880 109380 189120 109400
rect 189380 109380 189620 109400
rect 189880 109380 190120 109400
rect 190380 109380 190620 109400
rect 190880 109380 191120 109400
rect 191380 109380 191620 109400
rect 191880 109380 192120 109400
rect 192380 109380 192620 109400
rect 192880 109380 193120 109400
rect 193380 109380 193620 109400
rect 193880 109380 194120 109400
rect 194380 109380 194620 109400
rect 194880 109380 195120 109400
rect 195380 109380 195620 109400
rect 195880 109380 196120 109400
rect 196380 109380 196620 109400
rect 196880 109380 197120 109400
rect 197380 109380 197620 109400
rect 197880 109380 198120 109400
rect 198380 109380 198620 109400
rect 198880 109380 199120 109400
rect 199380 109380 199620 109400
rect 199880 109380 200120 109400
rect 200380 109380 200620 109400
rect 200880 109380 201120 109400
rect 201380 109380 201620 109400
rect 201880 109380 202120 109400
rect 202380 109380 202620 109400
rect 202880 109380 203120 109400
rect 203380 109380 203620 109400
rect 203880 109380 204120 109400
rect 204380 109380 204620 109400
rect 204880 109380 205120 109400
rect 205380 109380 205620 109400
rect 205880 109380 206120 109400
rect 206380 109380 206620 109400
rect 206880 109380 207120 109400
rect 207380 109380 207620 109400
rect 207880 109380 208120 109400
rect 208380 109380 208620 109400
rect 208880 109380 209120 109400
rect 209380 109380 209620 109400
rect 209880 109380 210120 109400
rect 210380 109380 210620 109400
rect 210880 109380 211120 109400
rect 211380 109380 211620 109400
rect 211880 109380 212120 109400
rect 212380 109380 212620 109400
rect 212880 109380 213120 109400
rect 213380 109380 213620 109400
rect 213880 109380 214120 109400
rect 214380 109380 214620 109400
rect 214880 109380 215120 109400
rect 215380 109380 215620 109400
rect 215880 109380 216120 109400
rect 216380 109380 216620 109400
rect 216880 109380 217120 109400
rect 217380 109380 217620 109400
rect 217880 109380 218120 109400
rect 218380 109380 218620 109400
rect 218880 109380 219120 109400
rect 219380 109380 219620 109400
rect 219880 109380 220120 109400
rect 220380 109380 220620 109400
rect 220880 109380 221120 109400
rect 221380 109380 221620 109400
rect 221880 109380 222120 109400
rect 222380 109380 222620 109400
rect 222880 109380 223120 109400
rect 223380 109380 223620 109400
rect 223880 109380 224120 109400
rect 224380 109380 224620 109400
rect 224880 109380 225120 109400
rect 225380 109380 225620 109400
rect 225880 109380 226120 109400
rect 226380 109380 226620 109400
rect 226880 109380 227120 109400
rect 227380 109380 227620 109400
rect 227880 109380 228120 109400
rect 228380 109380 228620 109400
rect 228880 109380 229120 109400
rect 229380 109380 229620 109400
rect 229880 109380 230120 109400
rect 230380 109380 230620 109400
rect 230880 109380 231120 109400
rect 231380 109380 231620 109400
rect 231880 109380 232000 109400
rect 178000 109120 178100 109380
rect 178400 109120 178600 109380
rect 178900 109120 179100 109380
rect 179400 109120 179600 109380
rect 179900 109120 180100 109380
rect 180400 109120 180600 109380
rect 180900 109120 181100 109380
rect 181400 109120 181600 109380
rect 181900 109120 182100 109380
rect 182400 109120 182600 109380
rect 182900 109120 183100 109380
rect 183400 109120 183600 109380
rect 183900 109120 184100 109380
rect 184400 109120 184600 109380
rect 184900 109120 185100 109380
rect 185400 109120 185600 109380
rect 185900 109120 186100 109380
rect 186400 109120 186600 109380
rect 186900 109120 187100 109380
rect 187400 109120 187600 109380
rect 187900 109120 188100 109380
rect 188400 109120 188600 109380
rect 188900 109120 189100 109380
rect 189400 109120 189600 109380
rect 189900 109120 190100 109380
rect 190400 109120 190600 109380
rect 190900 109120 191100 109380
rect 191400 109120 191600 109380
rect 191900 109120 192100 109380
rect 192400 109120 192600 109380
rect 192900 109120 193100 109380
rect 193400 109120 193600 109380
rect 193900 109120 194100 109380
rect 194400 109120 194600 109380
rect 194900 109120 195100 109380
rect 195400 109120 195600 109380
rect 195900 109120 196100 109380
rect 196400 109120 196600 109380
rect 196900 109120 197100 109380
rect 197400 109120 197600 109380
rect 197900 109120 198100 109380
rect 198400 109120 198600 109380
rect 198900 109120 199100 109380
rect 199400 109120 199600 109380
rect 199900 109120 200100 109380
rect 200400 109120 200600 109380
rect 200900 109120 201100 109380
rect 201400 109120 201600 109380
rect 201900 109120 202100 109380
rect 202400 109120 202600 109380
rect 202900 109120 203100 109380
rect 203400 109120 203600 109380
rect 203900 109120 204100 109380
rect 204400 109120 204600 109380
rect 204900 109120 205100 109380
rect 205400 109120 205600 109380
rect 205900 109120 206100 109380
rect 206400 109120 206600 109380
rect 206900 109120 207100 109380
rect 207400 109120 207600 109380
rect 207900 109120 208100 109380
rect 208400 109120 208600 109380
rect 208900 109120 209100 109380
rect 209400 109120 209600 109380
rect 209900 109120 210100 109380
rect 210400 109120 210600 109380
rect 210900 109120 211100 109380
rect 211400 109120 211600 109380
rect 211900 109120 212100 109380
rect 212400 109120 212600 109380
rect 212900 109120 213100 109380
rect 213400 109120 213600 109380
rect 213900 109120 214100 109380
rect 214400 109120 214600 109380
rect 214900 109120 215100 109380
rect 215400 109120 215600 109380
rect 215900 109120 216100 109380
rect 216400 109120 216600 109380
rect 216900 109120 217100 109380
rect 217400 109120 217600 109380
rect 217900 109120 218100 109380
rect 218400 109120 218600 109380
rect 218900 109120 219100 109380
rect 219400 109120 219600 109380
rect 219900 109120 220100 109380
rect 220400 109120 220600 109380
rect 220900 109120 221100 109380
rect 221400 109120 221600 109380
rect 221900 109120 222100 109380
rect 222400 109120 222600 109380
rect 222900 109120 223100 109380
rect 223400 109120 223600 109380
rect 223900 109120 224100 109380
rect 224400 109120 224600 109380
rect 224900 109120 225100 109380
rect 225400 109120 225600 109380
rect 225900 109120 226100 109380
rect 226400 109120 226600 109380
rect 226900 109120 227100 109380
rect 227400 109120 227600 109380
rect 227900 109120 228100 109380
rect 228400 109120 228600 109380
rect 228900 109120 229100 109380
rect 229400 109120 229600 109380
rect 229900 109120 230100 109380
rect 230400 109120 230600 109380
rect 230900 109120 231100 109380
rect 231400 109120 231600 109380
rect 231900 109120 232000 109380
rect 178000 109100 178120 109120
rect 178380 109100 178620 109120
rect 178880 109100 179120 109120
rect 179380 109100 179620 109120
rect 179880 109100 180120 109120
rect 180380 109100 180620 109120
rect 180880 109100 181120 109120
rect 181380 109100 181620 109120
rect 181880 109100 182120 109120
rect 182380 109100 182620 109120
rect 182880 109100 183120 109120
rect 183380 109100 183620 109120
rect 183880 109100 184120 109120
rect 184380 109100 184620 109120
rect 184880 109100 185120 109120
rect 185380 109100 185620 109120
rect 185880 109100 186120 109120
rect 186380 109100 186620 109120
rect 186880 109100 187120 109120
rect 187380 109100 187620 109120
rect 187880 109100 188120 109120
rect 188380 109100 188620 109120
rect 188880 109100 189120 109120
rect 189380 109100 189620 109120
rect 189880 109100 190120 109120
rect 190380 109100 190620 109120
rect 190880 109100 191120 109120
rect 191380 109100 191620 109120
rect 191880 109100 192120 109120
rect 192380 109100 192620 109120
rect 192880 109100 193120 109120
rect 193380 109100 193620 109120
rect 193880 109100 194120 109120
rect 194380 109100 194620 109120
rect 194880 109100 195120 109120
rect 195380 109100 195620 109120
rect 195880 109100 196120 109120
rect 196380 109100 196620 109120
rect 196880 109100 197120 109120
rect 197380 109100 197620 109120
rect 197880 109100 198120 109120
rect 198380 109100 198620 109120
rect 198880 109100 199120 109120
rect 199380 109100 199620 109120
rect 199880 109100 200120 109120
rect 200380 109100 200620 109120
rect 200880 109100 201120 109120
rect 201380 109100 201620 109120
rect 201880 109100 202120 109120
rect 202380 109100 202620 109120
rect 202880 109100 203120 109120
rect 203380 109100 203620 109120
rect 203880 109100 204120 109120
rect 204380 109100 204620 109120
rect 204880 109100 205120 109120
rect 205380 109100 205620 109120
rect 205880 109100 206120 109120
rect 206380 109100 206620 109120
rect 206880 109100 207120 109120
rect 207380 109100 207620 109120
rect 207880 109100 208120 109120
rect 208380 109100 208620 109120
rect 208880 109100 209120 109120
rect 209380 109100 209620 109120
rect 209880 109100 210120 109120
rect 210380 109100 210620 109120
rect 210880 109100 211120 109120
rect 211380 109100 211620 109120
rect 211880 109100 212120 109120
rect 212380 109100 212620 109120
rect 212880 109100 213120 109120
rect 213380 109100 213620 109120
rect 213880 109100 214120 109120
rect 214380 109100 214620 109120
rect 214880 109100 215120 109120
rect 215380 109100 215620 109120
rect 215880 109100 216120 109120
rect 216380 109100 216620 109120
rect 216880 109100 217120 109120
rect 217380 109100 217620 109120
rect 217880 109100 218120 109120
rect 218380 109100 218620 109120
rect 218880 109100 219120 109120
rect 219380 109100 219620 109120
rect 219880 109100 220120 109120
rect 220380 109100 220620 109120
rect 220880 109100 221120 109120
rect 221380 109100 221620 109120
rect 221880 109100 222120 109120
rect 222380 109100 222620 109120
rect 222880 109100 223120 109120
rect 223380 109100 223620 109120
rect 223880 109100 224120 109120
rect 224380 109100 224620 109120
rect 224880 109100 225120 109120
rect 225380 109100 225620 109120
rect 225880 109100 226120 109120
rect 226380 109100 226620 109120
rect 226880 109100 227120 109120
rect 227380 109100 227620 109120
rect 227880 109100 228120 109120
rect 228380 109100 228620 109120
rect 228880 109100 229120 109120
rect 229380 109100 229620 109120
rect 229880 109100 230120 109120
rect 230380 109100 230620 109120
rect 230880 109100 231120 109120
rect 231380 109100 231620 109120
rect 231880 109100 232000 109120
rect 178000 108900 232000 109100
rect 178000 108880 178120 108900
rect 178380 108880 178620 108900
rect 178880 108880 179120 108900
rect 179380 108880 179620 108900
rect 179880 108880 180120 108900
rect 180380 108880 180620 108900
rect 180880 108880 181120 108900
rect 181380 108880 181620 108900
rect 181880 108880 182120 108900
rect 182380 108880 182620 108900
rect 182880 108880 183120 108900
rect 183380 108880 183620 108900
rect 183880 108880 184120 108900
rect 184380 108880 184620 108900
rect 184880 108880 185120 108900
rect 185380 108880 185620 108900
rect 185880 108880 186120 108900
rect 186380 108880 186620 108900
rect 186880 108880 187120 108900
rect 187380 108880 187620 108900
rect 187880 108880 188120 108900
rect 188380 108880 188620 108900
rect 188880 108880 189120 108900
rect 189380 108880 189620 108900
rect 189880 108880 190120 108900
rect 190380 108880 190620 108900
rect 190880 108880 191120 108900
rect 191380 108880 191620 108900
rect 191880 108880 192120 108900
rect 192380 108880 192620 108900
rect 192880 108880 193120 108900
rect 193380 108880 193620 108900
rect 193880 108880 194120 108900
rect 194380 108880 194620 108900
rect 194880 108880 195120 108900
rect 195380 108880 195620 108900
rect 195880 108880 196120 108900
rect 196380 108880 196620 108900
rect 196880 108880 197120 108900
rect 197380 108880 197620 108900
rect 197880 108880 198120 108900
rect 198380 108880 198620 108900
rect 198880 108880 199120 108900
rect 199380 108880 199620 108900
rect 199880 108880 200120 108900
rect 200380 108880 200620 108900
rect 200880 108880 201120 108900
rect 201380 108880 201620 108900
rect 201880 108880 202120 108900
rect 202380 108880 202620 108900
rect 202880 108880 203120 108900
rect 203380 108880 203620 108900
rect 203880 108880 204120 108900
rect 204380 108880 204620 108900
rect 204880 108880 205120 108900
rect 205380 108880 205620 108900
rect 205880 108880 206120 108900
rect 206380 108880 206620 108900
rect 206880 108880 207120 108900
rect 207380 108880 207620 108900
rect 207880 108880 208120 108900
rect 208380 108880 208620 108900
rect 208880 108880 209120 108900
rect 209380 108880 209620 108900
rect 209880 108880 210120 108900
rect 210380 108880 210620 108900
rect 210880 108880 211120 108900
rect 211380 108880 211620 108900
rect 211880 108880 212120 108900
rect 212380 108880 212620 108900
rect 212880 108880 213120 108900
rect 213380 108880 213620 108900
rect 213880 108880 214120 108900
rect 214380 108880 214620 108900
rect 214880 108880 215120 108900
rect 215380 108880 215620 108900
rect 215880 108880 216120 108900
rect 216380 108880 216620 108900
rect 216880 108880 217120 108900
rect 217380 108880 217620 108900
rect 217880 108880 218120 108900
rect 218380 108880 218620 108900
rect 218880 108880 219120 108900
rect 219380 108880 219620 108900
rect 219880 108880 220120 108900
rect 220380 108880 220620 108900
rect 220880 108880 221120 108900
rect 221380 108880 221620 108900
rect 221880 108880 222120 108900
rect 222380 108880 222620 108900
rect 222880 108880 223120 108900
rect 223380 108880 223620 108900
rect 223880 108880 224120 108900
rect 224380 108880 224620 108900
rect 224880 108880 225120 108900
rect 225380 108880 225620 108900
rect 225880 108880 226120 108900
rect 226380 108880 226620 108900
rect 226880 108880 227120 108900
rect 227380 108880 227620 108900
rect 227880 108880 228120 108900
rect 228380 108880 228620 108900
rect 228880 108880 229120 108900
rect 229380 108880 229620 108900
rect 229880 108880 230120 108900
rect 230380 108880 230620 108900
rect 230880 108880 231120 108900
rect 231380 108880 231620 108900
rect 231880 108880 232000 108900
rect 178000 108620 178100 108880
rect 178400 108620 178600 108880
rect 178900 108620 179100 108880
rect 179400 108620 179600 108880
rect 179900 108620 180100 108880
rect 180400 108620 180600 108880
rect 180900 108620 181100 108880
rect 181400 108620 181600 108880
rect 181900 108620 182100 108880
rect 182400 108620 182600 108880
rect 182900 108620 183100 108880
rect 183400 108620 183600 108880
rect 183900 108620 184100 108880
rect 184400 108620 184600 108880
rect 184900 108620 185100 108880
rect 185400 108620 185600 108880
rect 185900 108620 186100 108880
rect 186400 108620 186600 108880
rect 186900 108620 187100 108880
rect 187400 108620 187600 108880
rect 187900 108620 188100 108880
rect 188400 108620 188600 108880
rect 188900 108620 189100 108880
rect 189400 108620 189600 108880
rect 189900 108620 190100 108880
rect 190400 108620 190600 108880
rect 190900 108620 191100 108880
rect 191400 108620 191600 108880
rect 191900 108620 192100 108880
rect 192400 108620 192600 108880
rect 192900 108620 193100 108880
rect 193400 108620 193600 108880
rect 193900 108620 194100 108880
rect 194400 108620 194600 108880
rect 194900 108620 195100 108880
rect 195400 108620 195600 108880
rect 195900 108620 196100 108880
rect 196400 108620 196600 108880
rect 196900 108620 197100 108880
rect 197400 108620 197600 108880
rect 197900 108620 198100 108880
rect 198400 108620 198600 108880
rect 198900 108620 199100 108880
rect 199400 108620 199600 108880
rect 199900 108620 200100 108880
rect 200400 108620 200600 108880
rect 200900 108620 201100 108880
rect 201400 108620 201600 108880
rect 201900 108620 202100 108880
rect 202400 108620 202600 108880
rect 202900 108620 203100 108880
rect 203400 108620 203600 108880
rect 203900 108620 204100 108880
rect 204400 108620 204600 108880
rect 204900 108620 205100 108880
rect 205400 108620 205600 108880
rect 205900 108620 206100 108880
rect 206400 108620 206600 108880
rect 206900 108620 207100 108880
rect 207400 108620 207600 108880
rect 207900 108620 208100 108880
rect 208400 108620 208600 108880
rect 208900 108620 209100 108880
rect 209400 108620 209600 108880
rect 209900 108620 210100 108880
rect 210400 108620 210600 108880
rect 210900 108620 211100 108880
rect 211400 108620 211600 108880
rect 211900 108620 212100 108880
rect 212400 108620 212600 108880
rect 212900 108620 213100 108880
rect 213400 108620 213600 108880
rect 213900 108620 214100 108880
rect 214400 108620 214600 108880
rect 214900 108620 215100 108880
rect 215400 108620 215600 108880
rect 215900 108620 216100 108880
rect 216400 108620 216600 108880
rect 216900 108620 217100 108880
rect 217400 108620 217600 108880
rect 217900 108620 218100 108880
rect 218400 108620 218600 108880
rect 218900 108620 219100 108880
rect 219400 108620 219600 108880
rect 219900 108620 220100 108880
rect 220400 108620 220600 108880
rect 220900 108620 221100 108880
rect 221400 108620 221600 108880
rect 221900 108620 222100 108880
rect 222400 108620 222600 108880
rect 222900 108620 223100 108880
rect 223400 108620 223600 108880
rect 223900 108620 224100 108880
rect 224400 108620 224600 108880
rect 224900 108620 225100 108880
rect 225400 108620 225600 108880
rect 225900 108620 226100 108880
rect 226400 108620 226600 108880
rect 226900 108620 227100 108880
rect 227400 108620 227600 108880
rect 227900 108620 228100 108880
rect 228400 108620 228600 108880
rect 228900 108620 229100 108880
rect 229400 108620 229600 108880
rect 229900 108620 230100 108880
rect 230400 108620 230600 108880
rect 230900 108620 231100 108880
rect 231400 108620 231600 108880
rect 231900 108620 232000 108880
rect 178000 108600 178120 108620
rect 178380 108600 178620 108620
rect 178880 108600 179120 108620
rect 179380 108600 179620 108620
rect 179880 108600 180120 108620
rect 180380 108600 180620 108620
rect 180880 108600 181120 108620
rect 181380 108600 181620 108620
rect 181880 108600 182120 108620
rect 182380 108600 182620 108620
rect 182880 108600 183120 108620
rect 183380 108600 183620 108620
rect 183880 108600 184120 108620
rect 184380 108600 184620 108620
rect 184880 108600 185120 108620
rect 185380 108600 185620 108620
rect 185880 108600 186120 108620
rect 186380 108600 186620 108620
rect 186880 108600 187120 108620
rect 187380 108600 187620 108620
rect 187880 108600 188120 108620
rect 188380 108600 188620 108620
rect 188880 108600 189120 108620
rect 189380 108600 189620 108620
rect 189880 108600 190120 108620
rect 190380 108600 190620 108620
rect 190880 108600 191120 108620
rect 191380 108600 191620 108620
rect 191880 108600 192120 108620
rect 192380 108600 192620 108620
rect 192880 108600 193120 108620
rect 193380 108600 193620 108620
rect 193880 108600 194120 108620
rect 194380 108600 194620 108620
rect 194880 108600 195120 108620
rect 195380 108600 195620 108620
rect 195880 108600 196120 108620
rect 196380 108600 196620 108620
rect 196880 108600 197120 108620
rect 197380 108600 197620 108620
rect 197880 108600 198120 108620
rect 198380 108600 198620 108620
rect 198880 108600 199120 108620
rect 199380 108600 199620 108620
rect 199880 108600 200120 108620
rect 200380 108600 200620 108620
rect 200880 108600 201120 108620
rect 201380 108600 201620 108620
rect 201880 108600 202120 108620
rect 202380 108600 202620 108620
rect 202880 108600 203120 108620
rect 203380 108600 203620 108620
rect 203880 108600 204120 108620
rect 204380 108600 204620 108620
rect 204880 108600 205120 108620
rect 205380 108600 205620 108620
rect 205880 108600 206120 108620
rect 206380 108600 206620 108620
rect 206880 108600 207120 108620
rect 207380 108600 207620 108620
rect 207880 108600 208120 108620
rect 208380 108600 208620 108620
rect 208880 108600 209120 108620
rect 209380 108600 209620 108620
rect 209880 108600 210120 108620
rect 210380 108600 210620 108620
rect 210880 108600 211120 108620
rect 211380 108600 211620 108620
rect 211880 108600 212120 108620
rect 212380 108600 212620 108620
rect 212880 108600 213120 108620
rect 213380 108600 213620 108620
rect 213880 108600 214120 108620
rect 214380 108600 214620 108620
rect 214880 108600 215120 108620
rect 215380 108600 215620 108620
rect 215880 108600 216120 108620
rect 216380 108600 216620 108620
rect 216880 108600 217120 108620
rect 217380 108600 217620 108620
rect 217880 108600 218120 108620
rect 218380 108600 218620 108620
rect 218880 108600 219120 108620
rect 219380 108600 219620 108620
rect 219880 108600 220120 108620
rect 220380 108600 220620 108620
rect 220880 108600 221120 108620
rect 221380 108600 221620 108620
rect 221880 108600 222120 108620
rect 222380 108600 222620 108620
rect 222880 108600 223120 108620
rect 223380 108600 223620 108620
rect 223880 108600 224120 108620
rect 224380 108600 224620 108620
rect 224880 108600 225120 108620
rect 225380 108600 225620 108620
rect 225880 108600 226120 108620
rect 226380 108600 226620 108620
rect 226880 108600 227120 108620
rect 227380 108600 227620 108620
rect 227880 108600 228120 108620
rect 228380 108600 228620 108620
rect 228880 108600 229120 108620
rect 229380 108600 229620 108620
rect 229880 108600 230120 108620
rect 230380 108600 230620 108620
rect 230880 108600 231120 108620
rect 231380 108600 231620 108620
rect 231880 108600 232000 108620
rect 178000 108400 232000 108600
rect 178000 108380 178120 108400
rect 178380 108380 178620 108400
rect 178880 108380 179120 108400
rect 179380 108380 179620 108400
rect 179880 108380 180120 108400
rect 180380 108380 180620 108400
rect 180880 108380 181120 108400
rect 181380 108380 181620 108400
rect 181880 108380 182120 108400
rect 182380 108380 182620 108400
rect 182880 108380 183120 108400
rect 183380 108380 183620 108400
rect 183880 108380 184120 108400
rect 184380 108380 184620 108400
rect 184880 108380 185120 108400
rect 185380 108380 185620 108400
rect 185880 108380 186120 108400
rect 186380 108380 186620 108400
rect 186880 108380 187120 108400
rect 187380 108380 187620 108400
rect 187880 108380 188120 108400
rect 188380 108380 188620 108400
rect 188880 108380 189120 108400
rect 189380 108380 189620 108400
rect 189880 108380 190120 108400
rect 190380 108380 190620 108400
rect 190880 108380 191120 108400
rect 191380 108380 191620 108400
rect 191880 108380 192120 108400
rect 192380 108380 192620 108400
rect 192880 108380 193120 108400
rect 193380 108380 193620 108400
rect 193880 108380 194120 108400
rect 194380 108380 194620 108400
rect 194880 108380 195120 108400
rect 195380 108380 195620 108400
rect 195880 108380 196120 108400
rect 196380 108380 196620 108400
rect 196880 108380 197120 108400
rect 197380 108380 197620 108400
rect 197880 108380 198120 108400
rect 198380 108380 198620 108400
rect 198880 108380 199120 108400
rect 199380 108380 199620 108400
rect 199880 108380 200120 108400
rect 200380 108380 200620 108400
rect 200880 108380 201120 108400
rect 201380 108380 201620 108400
rect 201880 108380 202120 108400
rect 202380 108380 202620 108400
rect 202880 108380 203120 108400
rect 203380 108380 203620 108400
rect 203880 108380 204120 108400
rect 204380 108380 204620 108400
rect 204880 108380 205120 108400
rect 205380 108380 205620 108400
rect 205880 108380 206120 108400
rect 206380 108380 206620 108400
rect 206880 108380 207120 108400
rect 207380 108380 207620 108400
rect 207880 108380 208120 108400
rect 208380 108380 208620 108400
rect 208880 108380 209120 108400
rect 209380 108380 209620 108400
rect 209880 108380 210120 108400
rect 210380 108380 210620 108400
rect 210880 108380 211120 108400
rect 211380 108380 211620 108400
rect 211880 108380 212120 108400
rect 212380 108380 212620 108400
rect 212880 108380 213120 108400
rect 213380 108380 213620 108400
rect 213880 108380 214120 108400
rect 214380 108380 214620 108400
rect 214880 108380 215120 108400
rect 215380 108380 215620 108400
rect 215880 108380 216120 108400
rect 216380 108380 216620 108400
rect 216880 108380 217120 108400
rect 217380 108380 217620 108400
rect 217880 108380 218120 108400
rect 218380 108380 218620 108400
rect 218880 108380 219120 108400
rect 219380 108380 219620 108400
rect 219880 108380 220120 108400
rect 220380 108380 220620 108400
rect 220880 108380 221120 108400
rect 221380 108380 221620 108400
rect 221880 108380 222120 108400
rect 222380 108380 222620 108400
rect 222880 108380 223120 108400
rect 223380 108380 223620 108400
rect 223880 108380 224120 108400
rect 224380 108380 224620 108400
rect 224880 108380 225120 108400
rect 225380 108380 225620 108400
rect 225880 108380 226120 108400
rect 226380 108380 226620 108400
rect 226880 108380 227120 108400
rect 227380 108380 227620 108400
rect 227880 108380 228120 108400
rect 228380 108380 228620 108400
rect 228880 108380 229120 108400
rect 229380 108380 229620 108400
rect 229880 108380 230120 108400
rect 230380 108380 230620 108400
rect 230880 108380 231120 108400
rect 231380 108380 231620 108400
rect 231880 108380 232000 108400
rect 178000 108120 178100 108380
rect 178400 108120 178600 108380
rect 178900 108120 179100 108380
rect 179400 108120 179600 108380
rect 179900 108120 180100 108380
rect 180400 108120 180600 108380
rect 180900 108120 181100 108380
rect 181400 108120 181600 108380
rect 181900 108120 182100 108380
rect 182400 108120 182600 108380
rect 182900 108120 183100 108380
rect 183400 108120 183600 108380
rect 183900 108120 184100 108380
rect 184400 108120 184600 108380
rect 184900 108120 185100 108380
rect 185400 108120 185600 108380
rect 185900 108120 186100 108380
rect 186400 108120 186600 108380
rect 186900 108120 187100 108380
rect 187400 108120 187600 108380
rect 187900 108120 188100 108380
rect 188400 108120 188600 108380
rect 188900 108120 189100 108380
rect 189400 108120 189600 108380
rect 189900 108120 190100 108380
rect 190400 108120 190600 108380
rect 190900 108120 191100 108380
rect 191400 108120 191600 108380
rect 191900 108120 192100 108380
rect 192400 108120 192600 108380
rect 192900 108120 193100 108380
rect 193400 108120 193600 108380
rect 193900 108120 194100 108380
rect 194400 108120 194600 108380
rect 194900 108120 195100 108380
rect 195400 108120 195600 108380
rect 195900 108120 196100 108380
rect 196400 108120 196600 108380
rect 196900 108120 197100 108380
rect 197400 108120 197600 108380
rect 197900 108120 198100 108380
rect 198400 108120 198600 108380
rect 198900 108120 199100 108380
rect 199400 108120 199600 108380
rect 199900 108120 200100 108380
rect 200400 108120 200600 108380
rect 200900 108120 201100 108380
rect 201400 108120 201600 108380
rect 201900 108120 202100 108380
rect 202400 108120 202600 108380
rect 202900 108120 203100 108380
rect 203400 108120 203600 108380
rect 203900 108120 204100 108380
rect 204400 108120 204600 108380
rect 204900 108120 205100 108380
rect 205400 108120 205600 108380
rect 205900 108120 206100 108380
rect 206400 108120 206600 108380
rect 206900 108120 207100 108380
rect 207400 108120 207600 108380
rect 207900 108120 208100 108380
rect 208400 108120 208600 108380
rect 208900 108120 209100 108380
rect 209400 108120 209600 108380
rect 209900 108120 210100 108380
rect 210400 108120 210600 108380
rect 210900 108120 211100 108380
rect 211400 108120 211600 108380
rect 211900 108120 212100 108380
rect 212400 108120 212600 108380
rect 212900 108120 213100 108380
rect 213400 108120 213600 108380
rect 213900 108120 214100 108380
rect 214400 108120 214600 108380
rect 214900 108120 215100 108380
rect 215400 108120 215600 108380
rect 215900 108120 216100 108380
rect 216400 108120 216600 108380
rect 216900 108120 217100 108380
rect 217400 108120 217600 108380
rect 217900 108120 218100 108380
rect 218400 108120 218600 108380
rect 218900 108120 219100 108380
rect 219400 108120 219600 108380
rect 219900 108120 220100 108380
rect 220400 108120 220600 108380
rect 220900 108120 221100 108380
rect 221400 108120 221600 108380
rect 221900 108120 222100 108380
rect 222400 108120 222600 108380
rect 222900 108120 223100 108380
rect 223400 108120 223600 108380
rect 223900 108120 224100 108380
rect 224400 108120 224600 108380
rect 224900 108120 225100 108380
rect 225400 108120 225600 108380
rect 225900 108120 226100 108380
rect 226400 108120 226600 108380
rect 226900 108120 227100 108380
rect 227400 108120 227600 108380
rect 227900 108120 228100 108380
rect 228400 108120 228600 108380
rect 228900 108120 229100 108380
rect 229400 108120 229600 108380
rect 229900 108120 230100 108380
rect 230400 108120 230600 108380
rect 230900 108120 231100 108380
rect 231400 108120 231600 108380
rect 231900 108120 232000 108380
rect 178000 108100 178120 108120
rect 178380 108100 178620 108120
rect 178880 108100 179120 108120
rect 179380 108100 179620 108120
rect 179880 108100 180120 108120
rect 180380 108100 180620 108120
rect 180880 108100 181120 108120
rect 181380 108100 181620 108120
rect 181880 108100 182120 108120
rect 182380 108100 182620 108120
rect 182880 108100 183120 108120
rect 183380 108100 183620 108120
rect 183880 108100 184120 108120
rect 184380 108100 184620 108120
rect 184880 108100 185120 108120
rect 185380 108100 185620 108120
rect 185880 108100 186120 108120
rect 186380 108100 186620 108120
rect 186880 108100 187120 108120
rect 187380 108100 187620 108120
rect 187880 108100 188120 108120
rect 188380 108100 188620 108120
rect 188880 108100 189120 108120
rect 189380 108100 189620 108120
rect 189880 108100 190120 108120
rect 190380 108100 190620 108120
rect 190880 108100 191120 108120
rect 191380 108100 191620 108120
rect 191880 108100 192120 108120
rect 192380 108100 192620 108120
rect 192880 108100 193120 108120
rect 193380 108100 193620 108120
rect 193880 108100 194120 108120
rect 194380 108100 194620 108120
rect 194880 108100 195120 108120
rect 195380 108100 195620 108120
rect 195880 108100 196120 108120
rect 196380 108100 196620 108120
rect 196880 108100 197120 108120
rect 197380 108100 197620 108120
rect 197880 108100 198120 108120
rect 198380 108100 198620 108120
rect 198880 108100 199120 108120
rect 199380 108100 199620 108120
rect 199880 108100 200120 108120
rect 200380 108100 200620 108120
rect 200880 108100 201120 108120
rect 201380 108100 201620 108120
rect 201880 108100 202120 108120
rect 202380 108100 202620 108120
rect 202880 108100 203120 108120
rect 203380 108100 203620 108120
rect 203880 108100 204120 108120
rect 204380 108100 204620 108120
rect 204880 108100 205120 108120
rect 205380 108100 205620 108120
rect 205880 108100 206120 108120
rect 206380 108100 206620 108120
rect 206880 108100 207120 108120
rect 207380 108100 207620 108120
rect 207880 108100 208120 108120
rect 208380 108100 208620 108120
rect 208880 108100 209120 108120
rect 209380 108100 209620 108120
rect 209880 108100 210120 108120
rect 210380 108100 210620 108120
rect 210880 108100 211120 108120
rect 211380 108100 211620 108120
rect 211880 108100 212120 108120
rect 212380 108100 212620 108120
rect 212880 108100 213120 108120
rect 213380 108100 213620 108120
rect 213880 108100 214120 108120
rect 214380 108100 214620 108120
rect 214880 108100 215120 108120
rect 215380 108100 215620 108120
rect 215880 108100 216120 108120
rect 216380 108100 216620 108120
rect 216880 108100 217120 108120
rect 217380 108100 217620 108120
rect 217880 108100 218120 108120
rect 218380 108100 218620 108120
rect 218880 108100 219120 108120
rect 219380 108100 219620 108120
rect 219880 108100 220120 108120
rect 220380 108100 220620 108120
rect 220880 108100 221120 108120
rect 221380 108100 221620 108120
rect 221880 108100 222120 108120
rect 222380 108100 222620 108120
rect 222880 108100 223120 108120
rect 223380 108100 223620 108120
rect 223880 108100 224120 108120
rect 224380 108100 224620 108120
rect 224880 108100 225120 108120
rect 225380 108100 225620 108120
rect 225880 108100 226120 108120
rect 226380 108100 226620 108120
rect 226880 108100 227120 108120
rect 227380 108100 227620 108120
rect 227880 108100 228120 108120
rect 228380 108100 228620 108120
rect 228880 108100 229120 108120
rect 229380 108100 229620 108120
rect 229880 108100 230120 108120
rect 230380 108100 230620 108120
rect 230880 108100 231120 108120
rect 231380 108100 231620 108120
rect 231880 108100 232000 108120
rect 178000 107900 232000 108100
rect 178000 107880 178120 107900
rect 178380 107880 178620 107900
rect 178880 107880 179120 107900
rect 179380 107880 179620 107900
rect 179880 107880 180120 107900
rect 180380 107880 180620 107900
rect 180880 107880 181120 107900
rect 181380 107880 181620 107900
rect 181880 107880 182120 107900
rect 182380 107880 182620 107900
rect 182880 107880 183120 107900
rect 183380 107880 183620 107900
rect 183880 107880 184120 107900
rect 184380 107880 184620 107900
rect 184880 107880 185120 107900
rect 185380 107880 185620 107900
rect 185880 107880 186120 107900
rect 186380 107880 186620 107900
rect 186880 107880 187120 107900
rect 187380 107880 187620 107900
rect 187880 107880 188120 107900
rect 188380 107880 188620 107900
rect 188880 107880 189120 107900
rect 189380 107880 189620 107900
rect 189880 107880 190120 107900
rect 190380 107880 190620 107900
rect 190880 107880 191120 107900
rect 191380 107880 191620 107900
rect 191880 107880 192120 107900
rect 192380 107880 192620 107900
rect 192880 107880 193120 107900
rect 193380 107880 193620 107900
rect 193880 107880 194120 107900
rect 194380 107880 194620 107900
rect 194880 107880 195120 107900
rect 195380 107880 195620 107900
rect 195880 107880 196120 107900
rect 196380 107880 196620 107900
rect 196880 107880 197120 107900
rect 197380 107880 197620 107900
rect 197880 107880 198120 107900
rect 198380 107880 198620 107900
rect 198880 107880 199120 107900
rect 199380 107880 199620 107900
rect 199880 107880 200120 107900
rect 200380 107880 200620 107900
rect 200880 107880 201120 107900
rect 201380 107880 201620 107900
rect 201880 107880 202120 107900
rect 202380 107880 202620 107900
rect 202880 107880 203120 107900
rect 203380 107880 203620 107900
rect 203880 107880 204120 107900
rect 204380 107880 204620 107900
rect 204880 107880 205120 107900
rect 205380 107880 205620 107900
rect 205880 107880 206120 107900
rect 206380 107880 206620 107900
rect 206880 107880 207120 107900
rect 207380 107880 207620 107900
rect 207880 107880 208120 107900
rect 208380 107880 208620 107900
rect 208880 107880 209120 107900
rect 209380 107880 209620 107900
rect 209880 107880 210120 107900
rect 210380 107880 210620 107900
rect 210880 107880 211120 107900
rect 211380 107880 211620 107900
rect 211880 107880 212120 107900
rect 212380 107880 212620 107900
rect 212880 107880 213120 107900
rect 213380 107880 213620 107900
rect 213880 107880 214120 107900
rect 214380 107880 214620 107900
rect 214880 107880 215120 107900
rect 215380 107880 215620 107900
rect 215880 107880 216120 107900
rect 216380 107880 216620 107900
rect 216880 107880 217120 107900
rect 217380 107880 217620 107900
rect 217880 107880 218120 107900
rect 218380 107880 218620 107900
rect 218880 107880 219120 107900
rect 219380 107880 219620 107900
rect 219880 107880 220120 107900
rect 220380 107880 220620 107900
rect 220880 107880 221120 107900
rect 221380 107880 221620 107900
rect 221880 107880 222120 107900
rect 222380 107880 222620 107900
rect 222880 107880 223120 107900
rect 223380 107880 223620 107900
rect 223880 107880 224120 107900
rect 224380 107880 224620 107900
rect 224880 107880 225120 107900
rect 225380 107880 225620 107900
rect 225880 107880 226120 107900
rect 226380 107880 226620 107900
rect 226880 107880 227120 107900
rect 227380 107880 227620 107900
rect 227880 107880 228120 107900
rect 228380 107880 228620 107900
rect 228880 107880 229120 107900
rect 229380 107880 229620 107900
rect 229880 107880 230120 107900
rect 230380 107880 230620 107900
rect 230880 107880 231120 107900
rect 231380 107880 231620 107900
rect 231880 107880 232000 107900
rect 178000 107620 178100 107880
rect 178400 107620 178600 107880
rect 178900 107620 179100 107880
rect 179400 107620 179600 107880
rect 179900 107620 180100 107880
rect 180400 107620 180600 107880
rect 180900 107620 181100 107880
rect 181400 107620 181600 107880
rect 181900 107620 182100 107880
rect 182400 107620 182600 107880
rect 182900 107620 183100 107880
rect 183400 107620 183600 107880
rect 183900 107620 184100 107880
rect 184400 107620 184600 107880
rect 184900 107620 185100 107880
rect 185400 107620 185600 107880
rect 185900 107620 186100 107880
rect 186400 107620 186600 107880
rect 186900 107620 187100 107880
rect 187400 107620 187600 107880
rect 187900 107620 188100 107880
rect 188400 107620 188600 107880
rect 188900 107620 189100 107880
rect 189400 107620 189600 107880
rect 189900 107620 190100 107880
rect 190400 107620 190600 107880
rect 190900 107620 191100 107880
rect 191400 107620 191600 107880
rect 191900 107620 192100 107880
rect 192400 107620 192600 107880
rect 192900 107620 193100 107880
rect 193400 107620 193600 107880
rect 193900 107620 194100 107880
rect 194400 107620 194600 107880
rect 194900 107620 195100 107880
rect 195400 107620 195600 107880
rect 195900 107620 196100 107880
rect 196400 107620 196600 107880
rect 196900 107620 197100 107880
rect 197400 107620 197600 107880
rect 197900 107620 198100 107880
rect 198400 107620 198600 107880
rect 198900 107620 199100 107880
rect 199400 107620 199600 107880
rect 199900 107620 200100 107880
rect 200400 107620 200600 107880
rect 200900 107620 201100 107880
rect 201400 107620 201600 107880
rect 201900 107620 202100 107880
rect 202400 107620 202600 107880
rect 202900 107620 203100 107880
rect 203400 107620 203600 107880
rect 203900 107620 204100 107880
rect 204400 107620 204600 107880
rect 204900 107620 205100 107880
rect 205400 107620 205600 107880
rect 205900 107620 206100 107880
rect 206400 107620 206600 107880
rect 206900 107620 207100 107880
rect 207400 107620 207600 107880
rect 207900 107620 208100 107880
rect 208400 107620 208600 107880
rect 208900 107620 209100 107880
rect 209400 107620 209600 107880
rect 209900 107620 210100 107880
rect 210400 107620 210600 107880
rect 210900 107620 211100 107880
rect 211400 107620 211600 107880
rect 211900 107620 212100 107880
rect 212400 107620 212600 107880
rect 212900 107620 213100 107880
rect 213400 107620 213600 107880
rect 213900 107620 214100 107880
rect 214400 107620 214600 107880
rect 214900 107620 215100 107880
rect 215400 107620 215600 107880
rect 215900 107620 216100 107880
rect 216400 107620 216600 107880
rect 216900 107620 217100 107880
rect 217400 107620 217600 107880
rect 217900 107620 218100 107880
rect 218400 107620 218600 107880
rect 218900 107620 219100 107880
rect 219400 107620 219600 107880
rect 219900 107620 220100 107880
rect 220400 107620 220600 107880
rect 220900 107620 221100 107880
rect 221400 107620 221600 107880
rect 221900 107620 222100 107880
rect 222400 107620 222600 107880
rect 222900 107620 223100 107880
rect 223400 107620 223600 107880
rect 223900 107620 224100 107880
rect 224400 107620 224600 107880
rect 224900 107620 225100 107880
rect 225400 107620 225600 107880
rect 225900 107620 226100 107880
rect 226400 107620 226600 107880
rect 226900 107620 227100 107880
rect 227400 107620 227600 107880
rect 227900 107620 228100 107880
rect 228400 107620 228600 107880
rect 228900 107620 229100 107880
rect 229400 107620 229600 107880
rect 229900 107620 230100 107880
rect 230400 107620 230600 107880
rect 230900 107620 231100 107880
rect 231400 107620 231600 107880
rect 231900 107620 232000 107880
rect 178000 107600 178120 107620
rect 178380 107600 178620 107620
rect 178880 107600 179120 107620
rect 179380 107600 179620 107620
rect 179880 107600 180120 107620
rect 180380 107600 180620 107620
rect 180880 107600 181120 107620
rect 181380 107600 181620 107620
rect 181880 107600 182120 107620
rect 182380 107600 182620 107620
rect 182880 107600 183120 107620
rect 183380 107600 183620 107620
rect 183880 107600 184120 107620
rect 184380 107600 184620 107620
rect 184880 107600 185120 107620
rect 185380 107600 185620 107620
rect 185880 107600 186120 107620
rect 186380 107600 186620 107620
rect 186880 107600 187120 107620
rect 187380 107600 187620 107620
rect 187880 107600 188120 107620
rect 188380 107600 188620 107620
rect 188880 107600 189120 107620
rect 189380 107600 189620 107620
rect 189880 107600 190120 107620
rect 190380 107600 190620 107620
rect 190880 107600 191120 107620
rect 191380 107600 191620 107620
rect 191880 107600 192120 107620
rect 192380 107600 192620 107620
rect 192880 107600 193120 107620
rect 193380 107600 193620 107620
rect 193880 107600 194120 107620
rect 194380 107600 194620 107620
rect 194880 107600 195120 107620
rect 195380 107600 195620 107620
rect 195880 107600 196120 107620
rect 196380 107600 196620 107620
rect 196880 107600 197120 107620
rect 197380 107600 197620 107620
rect 197880 107600 198120 107620
rect 198380 107600 198620 107620
rect 198880 107600 199120 107620
rect 199380 107600 199620 107620
rect 199880 107600 200120 107620
rect 200380 107600 200620 107620
rect 200880 107600 201120 107620
rect 201380 107600 201620 107620
rect 201880 107600 202120 107620
rect 202380 107600 202620 107620
rect 202880 107600 203120 107620
rect 203380 107600 203620 107620
rect 203880 107600 204120 107620
rect 204380 107600 204620 107620
rect 204880 107600 205120 107620
rect 205380 107600 205620 107620
rect 205880 107600 206120 107620
rect 206380 107600 206620 107620
rect 206880 107600 207120 107620
rect 207380 107600 207620 107620
rect 207880 107600 208120 107620
rect 208380 107600 208620 107620
rect 208880 107600 209120 107620
rect 209380 107600 209620 107620
rect 209880 107600 210120 107620
rect 210380 107600 210620 107620
rect 210880 107600 211120 107620
rect 211380 107600 211620 107620
rect 211880 107600 212120 107620
rect 212380 107600 212620 107620
rect 212880 107600 213120 107620
rect 213380 107600 213620 107620
rect 213880 107600 214120 107620
rect 214380 107600 214620 107620
rect 214880 107600 215120 107620
rect 215380 107600 215620 107620
rect 215880 107600 216120 107620
rect 216380 107600 216620 107620
rect 216880 107600 217120 107620
rect 217380 107600 217620 107620
rect 217880 107600 218120 107620
rect 218380 107600 218620 107620
rect 218880 107600 219120 107620
rect 219380 107600 219620 107620
rect 219880 107600 220120 107620
rect 220380 107600 220620 107620
rect 220880 107600 221120 107620
rect 221380 107600 221620 107620
rect 221880 107600 222120 107620
rect 222380 107600 222620 107620
rect 222880 107600 223120 107620
rect 223380 107600 223620 107620
rect 223880 107600 224120 107620
rect 224380 107600 224620 107620
rect 224880 107600 225120 107620
rect 225380 107600 225620 107620
rect 225880 107600 226120 107620
rect 226380 107600 226620 107620
rect 226880 107600 227120 107620
rect 227380 107600 227620 107620
rect 227880 107600 228120 107620
rect 228380 107600 228620 107620
rect 228880 107600 229120 107620
rect 229380 107600 229620 107620
rect 229880 107600 230120 107620
rect 230380 107600 230620 107620
rect 230880 107600 231120 107620
rect 231380 107600 231620 107620
rect 231880 107600 232000 107620
rect 178000 107400 232000 107600
rect 178000 107380 178120 107400
rect 178380 107380 178620 107400
rect 178880 107380 179120 107400
rect 179380 107380 179620 107400
rect 179880 107380 180120 107400
rect 180380 107380 180620 107400
rect 180880 107380 181120 107400
rect 181380 107380 181620 107400
rect 181880 107380 182120 107400
rect 182380 107380 182620 107400
rect 182880 107380 183120 107400
rect 183380 107380 183620 107400
rect 183880 107380 184120 107400
rect 184380 107380 184620 107400
rect 184880 107380 185120 107400
rect 185380 107380 185620 107400
rect 185880 107380 186120 107400
rect 186380 107380 186620 107400
rect 186880 107380 187120 107400
rect 187380 107380 187620 107400
rect 187880 107380 188120 107400
rect 188380 107380 188620 107400
rect 188880 107380 189120 107400
rect 189380 107380 189620 107400
rect 189880 107380 190120 107400
rect 190380 107380 190620 107400
rect 190880 107380 191120 107400
rect 191380 107380 191620 107400
rect 191880 107380 192120 107400
rect 192380 107380 192620 107400
rect 192880 107380 193120 107400
rect 193380 107380 193620 107400
rect 193880 107380 194120 107400
rect 194380 107380 194620 107400
rect 194880 107380 195120 107400
rect 195380 107380 195620 107400
rect 195880 107380 196120 107400
rect 196380 107380 196620 107400
rect 196880 107380 197120 107400
rect 197380 107380 197620 107400
rect 197880 107380 198120 107400
rect 198380 107380 198620 107400
rect 198880 107380 199120 107400
rect 199380 107380 199620 107400
rect 199880 107380 200120 107400
rect 200380 107380 200620 107400
rect 200880 107380 201120 107400
rect 201380 107380 201620 107400
rect 201880 107380 202120 107400
rect 202380 107380 202620 107400
rect 202880 107380 203120 107400
rect 203380 107380 203620 107400
rect 203880 107380 204120 107400
rect 204380 107380 204620 107400
rect 204880 107380 205120 107400
rect 205380 107380 205620 107400
rect 205880 107380 206120 107400
rect 206380 107380 206620 107400
rect 206880 107380 207120 107400
rect 207380 107380 207620 107400
rect 207880 107380 208120 107400
rect 208380 107380 208620 107400
rect 208880 107380 209120 107400
rect 209380 107380 209620 107400
rect 209880 107380 210120 107400
rect 210380 107380 210620 107400
rect 210880 107380 211120 107400
rect 211380 107380 211620 107400
rect 211880 107380 212120 107400
rect 212380 107380 212620 107400
rect 212880 107380 213120 107400
rect 213380 107380 213620 107400
rect 213880 107380 214120 107400
rect 214380 107380 214620 107400
rect 214880 107380 215120 107400
rect 215380 107380 215620 107400
rect 215880 107380 216120 107400
rect 216380 107380 216620 107400
rect 216880 107380 217120 107400
rect 217380 107380 217620 107400
rect 217880 107380 218120 107400
rect 218380 107380 218620 107400
rect 218880 107380 219120 107400
rect 219380 107380 219620 107400
rect 219880 107380 220120 107400
rect 220380 107380 220620 107400
rect 220880 107380 221120 107400
rect 221380 107380 221620 107400
rect 221880 107380 222120 107400
rect 222380 107380 222620 107400
rect 222880 107380 223120 107400
rect 223380 107380 223620 107400
rect 223880 107380 224120 107400
rect 224380 107380 224620 107400
rect 224880 107380 225120 107400
rect 225380 107380 225620 107400
rect 225880 107380 226120 107400
rect 226380 107380 226620 107400
rect 226880 107380 227120 107400
rect 227380 107380 227620 107400
rect 227880 107380 228120 107400
rect 228380 107380 228620 107400
rect 228880 107380 229120 107400
rect 229380 107380 229620 107400
rect 229880 107380 230120 107400
rect 230380 107380 230620 107400
rect 230880 107380 231120 107400
rect 231380 107380 231620 107400
rect 231880 107380 232000 107400
rect 178000 107120 178100 107380
rect 178400 107120 178600 107380
rect 178900 107120 179100 107380
rect 179400 107120 179600 107380
rect 179900 107120 180100 107380
rect 180400 107120 180600 107380
rect 180900 107120 181100 107380
rect 181400 107120 181600 107380
rect 181900 107120 182100 107380
rect 182400 107120 182600 107380
rect 182900 107120 183100 107380
rect 183400 107120 183600 107380
rect 183900 107120 184100 107380
rect 184400 107120 184600 107380
rect 184900 107120 185100 107380
rect 185400 107120 185600 107380
rect 185900 107120 186100 107380
rect 186400 107120 186600 107380
rect 186900 107120 187100 107380
rect 187400 107120 187600 107380
rect 187900 107120 188100 107380
rect 188400 107120 188600 107380
rect 188900 107120 189100 107380
rect 189400 107120 189600 107380
rect 189900 107120 190100 107380
rect 190400 107120 190600 107380
rect 190900 107120 191100 107380
rect 191400 107120 191600 107380
rect 191900 107120 192100 107380
rect 192400 107120 192600 107380
rect 192900 107120 193100 107380
rect 193400 107120 193600 107380
rect 193900 107120 194100 107380
rect 194400 107120 194600 107380
rect 194900 107120 195100 107380
rect 195400 107120 195600 107380
rect 195900 107120 196100 107380
rect 196400 107120 196600 107380
rect 196900 107120 197100 107380
rect 197400 107120 197600 107380
rect 197900 107120 198100 107380
rect 198400 107120 198600 107380
rect 198900 107120 199100 107380
rect 199400 107120 199600 107380
rect 199900 107120 200100 107380
rect 200400 107120 200600 107380
rect 200900 107120 201100 107380
rect 201400 107120 201600 107380
rect 201900 107120 202100 107380
rect 202400 107120 202600 107380
rect 202900 107120 203100 107380
rect 203400 107120 203600 107380
rect 203900 107120 204100 107380
rect 204400 107120 204600 107380
rect 204900 107120 205100 107380
rect 205400 107120 205600 107380
rect 205900 107120 206100 107380
rect 206400 107120 206600 107380
rect 206900 107120 207100 107380
rect 207400 107120 207600 107380
rect 207900 107120 208100 107380
rect 208400 107120 208600 107380
rect 208900 107120 209100 107380
rect 209400 107120 209600 107380
rect 209900 107120 210100 107380
rect 210400 107120 210600 107380
rect 210900 107120 211100 107380
rect 211400 107120 211600 107380
rect 211900 107120 212100 107380
rect 212400 107120 212600 107380
rect 212900 107120 213100 107380
rect 213400 107120 213600 107380
rect 213900 107120 214100 107380
rect 214400 107120 214600 107380
rect 214900 107120 215100 107380
rect 215400 107120 215600 107380
rect 215900 107120 216100 107380
rect 216400 107120 216600 107380
rect 216900 107120 217100 107380
rect 217400 107120 217600 107380
rect 217900 107120 218100 107380
rect 218400 107120 218600 107380
rect 218900 107120 219100 107380
rect 219400 107120 219600 107380
rect 219900 107120 220100 107380
rect 220400 107120 220600 107380
rect 220900 107120 221100 107380
rect 221400 107120 221600 107380
rect 221900 107120 222100 107380
rect 222400 107120 222600 107380
rect 222900 107120 223100 107380
rect 223400 107120 223600 107380
rect 223900 107120 224100 107380
rect 224400 107120 224600 107380
rect 224900 107120 225100 107380
rect 225400 107120 225600 107380
rect 225900 107120 226100 107380
rect 226400 107120 226600 107380
rect 226900 107120 227100 107380
rect 227400 107120 227600 107380
rect 227900 107120 228100 107380
rect 228400 107120 228600 107380
rect 228900 107120 229100 107380
rect 229400 107120 229600 107380
rect 229900 107120 230100 107380
rect 230400 107120 230600 107380
rect 230900 107120 231100 107380
rect 231400 107120 231600 107380
rect 231900 107120 232000 107380
rect 178000 107100 178120 107120
rect 178380 107100 178620 107120
rect 178880 107100 179120 107120
rect 179380 107100 179620 107120
rect 179880 107100 180120 107120
rect 180380 107100 180620 107120
rect 180880 107100 181120 107120
rect 181380 107100 181620 107120
rect 181880 107100 182120 107120
rect 182380 107100 182620 107120
rect 182880 107100 183120 107120
rect 183380 107100 183620 107120
rect 183880 107100 184120 107120
rect 184380 107100 184620 107120
rect 184880 107100 185120 107120
rect 185380 107100 185620 107120
rect 185880 107100 186120 107120
rect 186380 107100 186620 107120
rect 186880 107100 187120 107120
rect 187380 107100 187620 107120
rect 187880 107100 188120 107120
rect 188380 107100 188620 107120
rect 188880 107100 189120 107120
rect 189380 107100 189620 107120
rect 189880 107100 190120 107120
rect 190380 107100 190620 107120
rect 190880 107100 191120 107120
rect 191380 107100 191620 107120
rect 191880 107100 192120 107120
rect 192380 107100 192620 107120
rect 192880 107100 193120 107120
rect 193380 107100 193620 107120
rect 193880 107100 194120 107120
rect 194380 107100 194620 107120
rect 194880 107100 195120 107120
rect 195380 107100 195620 107120
rect 195880 107100 196120 107120
rect 196380 107100 196620 107120
rect 196880 107100 197120 107120
rect 197380 107100 197620 107120
rect 197880 107100 198120 107120
rect 198380 107100 198620 107120
rect 198880 107100 199120 107120
rect 199380 107100 199620 107120
rect 199880 107100 200120 107120
rect 200380 107100 200620 107120
rect 200880 107100 201120 107120
rect 201380 107100 201620 107120
rect 201880 107100 202120 107120
rect 202380 107100 202620 107120
rect 202880 107100 203120 107120
rect 203380 107100 203620 107120
rect 203880 107100 204120 107120
rect 204380 107100 204620 107120
rect 204880 107100 205120 107120
rect 205380 107100 205620 107120
rect 205880 107100 206120 107120
rect 206380 107100 206620 107120
rect 206880 107100 207120 107120
rect 207380 107100 207620 107120
rect 207880 107100 208120 107120
rect 208380 107100 208620 107120
rect 208880 107100 209120 107120
rect 209380 107100 209620 107120
rect 209880 107100 210120 107120
rect 210380 107100 210620 107120
rect 210880 107100 211120 107120
rect 211380 107100 211620 107120
rect 211880 107100 212120 107120
rect 212380 107100 212620 107120
rect 212880 107100 213120 107120
rect 213380 107100 213620 107120
rect 213880 107100 214120 107120
rect 214380 107100 214620 107120
rect 214880 107100 215120 107120
rect 215380 107100 215620 107120
rect 215880 107100 216120 107120
rect 216380 107100 216620 107120
rect 216880 107100 217120 107120
rect 217380 107100 217620 107120
rect 217880 107100 218120 107120
rect 218380 107100 218620 107120
rect 218880 107100 219120 107120
rect 219380 107100 219620 107120
rect 219880 107100 220120 107120
rect 220380 107100 220620 107120
rect 220880 107100 221120 107120
rect 221380 107100 221620 107120
rect 221880 107100 222120 107120
rect 222380 107100 222620 107120
rect 222880 107100 223120 107120
rect 223380 107100 223620 107120
rect 223880 107100 224120 107120
rect 224380 107100 224620 107120
rect 224880 107100 225120 107120
rect 225380 107100 225620 107120
rect 225880 107100 226120 107120
rect 226380 107100 226620 107120
rect 226880 107100 227120 107120
rect 227380 107100 227620 107120
rect 227880 107100 228120 107120
rect 228380 107100 228620 107120
rect 228880 107100 229120 107120
rect 229380 107100 229620 107120
rect 229880 107100 230120 107120
rect 230380 107100 230620 107120
rect 230880 107100 231120 107120
rect 231380 107100 231620 107120
rect 231880 107100 232000 107120
rect 178000 106900 232000 107100
rect 178000 106880 178120 106900
rect 178380 106880 178620 106900
rect 178880 106880 179120 106900
rect 179380 106880 179620 106900
rect 179880 106880 180120 106900
rect 180380 106880 180620 106900
rect 180880 106880 181120 106900
rect 181380 106880 181620 106900
rect 181880 106880 182120 106900
rect 182380 106880 182620 106900
rect 182880 106880 183120 106900
rect 183380 106880 183620 106900
rect 183880 106880 184120 106900
rect 184380 106880 184620 106900
rect 184880 106880 185120 106900
rect 185380 106880 185620 106900
rect 185880 106880 186120 106900
rect 186380 106880 186620 106900
rect 186880 106880 187120 106900
rect 187380 106880 187620 106900
rect 187880 106880 188120 106900
rect 188380 106880 188620 106900
rect 188880 106880 189120 106900
rect 189380 106880 189620 106900
rect 189880 106880 190120 106900
rect 190380 106880 190620 106900
rect 190880 106880 191120 106900
rect 191380 106880 191620 106900
rect 191880 106880 192120 106900
rect 192380 106880 192620 106900
rect 192880 106880 193120 106900
rect 193380 106880 193620 106900
rect 193880 106880 194120 106900
rect 194380 106880 194620 106900
rect 194880 106880 195120 106900
rect 195380 106880 195620 106900
rect 195880 106880 196120 106900
rect 196380 106880 196620 106900
rect 196880 106880 197120 106900
rect 197380 106880 197620 106900
rect 197880 106880 198120 106900
rect 198380 106880 198620 106900
rect 198880 106880 199120 106900
rect 199380 106880 199620 106900
rect 199880 106880 200120 106900
rect 200380 106880 200620 106900
rect 200880 106880 201120 106900
rect 201380 106880 201620 106900
rect 201880 106880 202120 106900
rect 202380 106880 202620 106900
rect 202880 106880 203120 106900
rect 203380 106880 203620 106900
rect 203880 106880 204120 106900
rect 204380 106880 204620 106900
rect 204880 106880 205120 106900
rect 205380 106880 205620 106900
rect 205880 106880 206120 106900
rect 206380 106880 206620 106900
rect 206880 106880 207120 106900
rect 207380 106880 207620 106900
rect 207880 106880 208120 106900
rect 208380 106880 208620 106900
rect 208880 106880 209120 106900
rect 209380 106880 209620 106900
rect 209880 106880 210120 106900
rect 210380 106880 210620 106900
rect 210880 106880 211120 106900
rect 211380 106880 211620 106900
rect 211880 106880 212120 106900
rect 212380 106880 212620 106900
rect 212880 106880 213120 106900
rect 213380 106880 213620 106900
rect 213880 106880 214120 106900
rect 214380 106880 214620 106900
rect 214880 106880 215120 106900
rect 215380 106880 215620 106900
rect 215880 106880 216120 106900
rect 216380 106880 216620 106900
rect 216880 106880 217120 106900
rect 217380 106880 217620 106900
rect 217880 106880 218120 106900
rect 218380 106880 218620 106900
rect 218880 106880 219120 106900
rect 219380 106880 219620 106900
rect 219880 106880 220120 106900
rect 220380 106880 220620 106900
rect 220880 106880 221120 106900
rect 221380 106880 221620 106900
rect 221880 106880 222120 106900
rect 222380 106880 222620 106900
rect 222880 106880 223120 106900
rect 223380 106880 223620 106900
rect 223880 106880 224120 106900
rect 224380 106880 224620 106900
rect 224880 106880 225120 106900
rect 225380 106880 225620 106900
rect 225880 106880 226120 106900
rect 226380 106880 226620 106900
rect 226880 106880 227120 106900
rect 227380 106880 227620 106900
rect 227880 106880 228120 106900
rect 228380 106880 228620 106900
rect 228880 106880 229120 106900
rect 229380 106880 229620 106900
rect 229880 106880 230120 106900
rect 230380 106880 230620 106900
rect 230880 106880 231120 106900
rect 231380 106880 231620 106900
rect 231880 106880 232000 106900
rect 178000 106620 178100 106880
rect 178400 106620 178600 106880
rect 178900 106620 179100 106880
rect 179400 106620 179600 106880
rect 179900 106620 180100 106880
rect 180400 106620 180600 106880
rect 180900 106620 181100 106880
rect 181400 106620 181600 106880
rect 181900 106620 182100 106880
rect 182400 106620 182600 106880
rect 182900 106620 183100 106880
rect 183400 106620 183600 106880
rect 183900 106620 184100 106880
rect 184400 106620 184600 106880
rect 184900 106620 185100 106880
rect 185400 106620 185600 106880
rect 185900 106620 186100 106880
rect 186400 106620 186600 106880
rect 186900 106620 187100 106880
rect 187400 106620 187600 106880
rect 187900 106620 188100 106880
rect 188400 106620 188600 106880
rect 188900 106620 189100 106880
rect 189400 106620 189600 106880
rect 189900 106620 190100 106880
rect 190400 106620 190600 106880
rect 190900 106620 191100 106880
rect 191400 106620 191600 106880
rect 191900 106620 192100 106880
rect 192400 106620 192600 106880
rect 192900 106620 193100 106880
rect 193400 106620 193600 106880
rect 193900 106620 194100 106880
rect 194400 106620 194600 106880
rect 194900 106620 195100 106880
rect 195400 106620 195600 106880
rect 195900 106620 196100 106880
rect 196400 106620 196600 106880
rect 196900 106620 197100 106880
rect 197400 106620 197600 106880
rect 197900 106620 198100 106880
rect 198400 106620 198600 106880
rect 198900 106620 199100 106880
rect 199400 106620 199600 106880
rect 199900 106620 200100 106880
rect 200400 106620 200600 106880
rect 200900 106620 201100 106880
rect 201400 106620 201600 106880
rect 201900 106620 202100 106880
rect 202400 106620 202600 106880
rect 202900 106620 203100 106880
rect 203400 106620 203600 106880
rect 203900 106620 204100 106880
rect 204400 106620 204600 106880
rect 204900 106620 205100 106880
rect 205400 106620 205600 106880
rect 205900 106620 206100 106880
rect 206400 106620 206600 106880
rect 206900 106620 207100 106880
rect 207400 106620 207600 106880
rect 207900 106620 208100 106880
rect 208400 106620 208600 106880
rect 208900 106620 209100 106880
rect 209400 106620 209600 106880
rect 209900 106620 210100 106880
rect 210400 106620 210600 106880
rect 210900 106620 211100 106880
rect 211400 106620 211600 106880
rect 211900 106620 212100 106880
rect 212400 106620 212600 106880
rect 212900 106620 213100 106880
rect 213400 106620 213600 106880
rect 213900 106620 214100 106880
rect 214400 106620 214600 106880
rect 214900 106620 215100 106880
rect 215400 106620 215600 106880
rect 215900 106620 216100 106880
rect 216400 106620 216600 106880
rect 216900 106620 217100 106880
rect 217400 106620 217600 106880
rect 217900 106620 218100 106880
rect 218400 106620 218600 106880
rect 218900 106620 219100 106880
rect 219400 106620 219600 106880
rect 219900 106620 220100 106880
rect 220400 106620 220600 106880
rect 220900 106620 221100 106880
rect 221400 106620 221600 106880
rect 221900 106620 222100 106880
rect 222400 106620 222600 106880
rect 222900 106620 223100 106880
rect 223400 106620 223600 106880
rect 223900 106620 224100 106880
rect 224400 106620 224600 106880
rect 224900 106620 225100 106880
rect 225400 106620 225600 106880
rect 225900 106620 226100 106880
rect 226400 106620 226600 106880
rect 226900 106620 227100 106880
rect 227400 106620 227600 106880
rect 227900 106620 228100 106880
rect 228400 106620 228600 106880
rect 228900 106620 229100 106880
rect 229400 106620 229600 106880
rect 229900 106620 230100 106880
rect 230400 106620 230600 106880
rect 230900 106620 231100 106880
rect 231400 106620 231600 106880
rect 231900 106620 232000 106880
rect 178000 106600 178120 106620
rect 178380 106600 178620 106620
rect 178880 106600 179120 106620
rect 179380 106600 179620 106620
rect 179880 106600 180120 106620
rect 180380 106600 180620 106620
rect 180880 106600 181120 106620
rect 181380 106600 181620 106620
rect 181880 106600 182120 106620
rect 182380 106600 182620 106620
rect 182880 106600 183120 106620
rect 183380 106600 183620 106620
rect 183880 106600 184120 106620
rect 184380 106600 184620 106620
rect 184880 106600 185120 106620
rect 185380 106600 185620 106620
rect 185880 106600 186120 106620
rect 186380 106600 186620 106620
rect 186880 106600 187120 106620
rect 187380 106600 187620 106620
rect 187880 106600 188120 106620
rect 188380 106600 188620 106620
rect 188880 106600 189120 106620
rect 189380 106600 189620 106620
rect 189880 106600 190120 106620
rect 190380 106600 190620 106620
rect 190880 106600 191120 106620
rect 191380 106600 191620 106620
rect 191880 106600 192120 106620
rect 192380 106600 192620 106620
rect 192880 106600 193120 106620
rect 193380 106600 193620 106620
rect 193880 106600 194120 106620
rect 194380 106600 194620 106620
rect 194880 106600 195120 106620
rect 195380 106600 195620 106620
rect 195880 106600 196120 106620
rect 196380 106600 196620 106620
rect 196880 106600 197120 106620
rect 197380 106600 197620 106620
rect 197880 106600 198120 106620
rect 198380 106600 198620 106620
rect 198880 106600 199120 106620
rect 199380 106600 199620 106620
rect 199880 106600 200120 106620
rect 200380 106600 200620 106620
rect 200880 106600 201120 106620
rect 201380 106600 201620 106620
rect 201880 106600 202120 106620
rect 202380 106600 202620 106620
rect 202880 106600 203120 106620
rect 203380 106600 203620 106620
rect 203880 106600 204120 106620
rect 204380 106600 204620 106620
rect 204880 106600 205120 106620
rect 205380 106600 205620 106620
rect 205880 106600 206120 106620
rect 206380 106600 206620 106620
rect 206880 106600 207120 106620
rect 207380 106600 207620 106620
rect 207880 106600 208120 106620
rect 208380 106600 208620 106620
rect 208880 106600 209120 106620
rect 209380 106600 209620 106620
rect 209880 106600 210120 106620
rect 210380 106600 210620 106620
rect 210880 106600 211120 106620
rect 211380 106600 211620 106620
rect 211880 106600 212120 106620
rect 212380 106600 212620 106620
rect 212880 106600 213120 106620
rect 213380 106600 213620 106620
rect 213880 106600 214120 106620
rect 214380 106600 214620 106620
rect 214880 106600 215120 106620
rect 215380 106600 215620 106620
rect 215880 106600 216120 106620
rect 216380 106600 216620 106620
rect 216880 106600 217120 106620
rect 217380 106600 217620 106620
rect 217880 106600 218120 106620
rect 218380 106600 218620 106620
rect 218880 106600 219120 106620
rect 219380 106600 219620 106620
rect 219880 106600 220120 106620
rect 220380 106600 220620 106620
rect 220880 106600 221120 106620
rect 221380 106600 221620 106620
rect 221880 106600 222120 106620
rect 222380 106600 222620 106620
rect 222880 106600 223120 106620
rect 223380 106600 223620 106620
rect 223880 106600 224120 106620
rect 224380 106600 224620 106620
rect 224880 106600 225120 106620
rect 225380 106600 225620 106620
rect 225880 106600 226120 106620
rect 226380 106600 226620 106620
rect 226880 106600 227120 106620
rect 227380 106600 227620 106620
rect 227880 106600 228120 106620
rect 228380 106600 228620 106620
rect 228880 106600 229120 106620
rect 229380 106600 229620 106620
rect 229880 106600 230120 106620
rect 230380 106600 230620 106620
rect 230880 106600 231120 106620
rect 231380 106600 231620 106620
rect 231880 106600 232000 106620
rect 178000 106400 232000 106600
rect 178000 106380 178120 106400
rect 178380 106380 178620 106400
rect 178880 106380 179120 106400
rect 179380 106380 179620 106400
rect 179880 106380 180120 106400
rect 180380 106380 180620 106400
rect 180880 106380 181120 106400
rect 181380 106380 181620 106400
rect 181880 106380 182120 106400
rect 182380 106380 182620 106400
rect 182880 106380 183120 106400
rect 183380 106380 183620 106400
rect 183880 106380 184120 106400
rect 184380 106380 184620 106400
rect 184880 106380 185120 106400
rect 185380 106380 185620 106400
rect 185880 106380 186120 106400
rect 186380 106380 186620 106400
rect 186880 106380 187120 106400
rect 187380 106380 187620 106400
rect 187880 106380 188120 106400
rect 188380 106380 188620 106400
rect 188880 106380 189120 106400
rect 189380 106380 189620 106400
rect 189880 106380 190120 106400
rect 190380 106380 190620 106400
rect 190880 106380 191120 106400
rect 191380 106380 191620 106400
rect 191880 106380 192120 106400
rect 192380 106380 192620 106400
rect 192880 106380 193120 106400
rect 193380 106380 193620 106400
rect 193880 106380 194120 106400
rect 194380 106380 194620 106400
rect 194880 106380 195120 106400
rect 195380 106380 195620 106400
rect 195880 106380 196120 106400
rect 196380 106380 196620 106400
rect 196880 106380 197120 106400
rect 197380 106380 197620 106400
rect 197880 106380 198120 106400
rect 198380 106380 198620 106400
rect 198880 106380 199120 106400
rect 199380 106380 199620 106400
rect 199880 106380 200120 106400
rect 200380 106380 200620 106400
rect 200880 106380 201120 106400
rect 201380 106380 201620 106400
rect 201880 106380 202120 106400
rect 202380 106380 202620 106400
rect 202880 106380 203120 106400
rect 203380 106380 203620 106400
rect 203880 106380 204120 106400
rect 204380 106380 204620 106400
rect 204880 106380 205120 106400
rect 205380 106380 205620 106400
rect 205880 106380 206120 106400
rect 206380 106380 206620 106400
rect 206880 106380 207120 106400
rect 207380 106380 207620 106400
rect 207880 106380 208120 106400
rect 208380 106380 208620 106400
rect 208880 106380 209120 106400
rect 209380 106380 209620 106400
rect 209880 106380 210120 106400
rect 210380 106380 210620 106400
rect 210880 106380 211120 106400
rect 211380 106380 211620 106400
rect 211880 106380 212120 106400
rect 212380 106380 212620 106400
rect 212880 106380 213120 106400
rect 213380 106380 213620 106400
rect 213880 106380 214120 106400
rect 214380 106380 214620 106400
rect 214880 106380 215120 106400
rect 215380 106380 215620 106400
rect 215880 106380 216120 106400
rect 216380 106380 216620 106400
rect 216880 106380 217120 106400
rect 217380 106380 217620 106400
rect 217880 106380 218120 106400
rect 218380 106380 218620 106400
rect 218880 106380 219120 106400
rect 219380 106380 219620 106400
rect 219880 106380 220120 106400
rect 220380 106380 220620 106400
rect 220880 106380 221120 106400
rect 221380 106380 221620 106400
rect 221880 106380 222120 106400
rect 222380 106380 222620 106400
rect 222880 106380 223120 106400
rect 223380 106380 223620 106400
rect 223880 106380 224120 106400
rect 224380 106380 224620 106400
rect 224880 106380 225120 106400
rect 225380 106380 225620 106400
rect 225880 106380 226120 106400
rect 226380 106380 226620 106400
rect 226880 106380 227120 106400
rect 227380 106380 227620 106400
rect 227880 106380 228120 106400
rect 228380 106380 228620 106400
rect 228880 106380 229120 106400
rect 229380 106380 229620 106400
rect 229880 106380 230120 106400
rect 230380 106380 230620 106400
rect 230880 106380 231120 106400
rect 231380 106380 231620 106400
rect 231880 106380 232000 106400
rect 178000 106120 178100 106380
rect 178400 106120 178600 106380
rect 178900 106120 179100 106380
rect 179400 106120 179600 106380
rect 179900 106120 180100 106380
rect 180400 106120 180600 106380
rect 180900 106120 181100 106380
rect 181400 106120 181600 106380
rect 181900 106120 182100 106380
rect 182400 106120 182600 106380
rect 182900 106120 183100 106380
rect 183400 106120 183600 106380
rect 183900 106120 184100 106380
rect 184400 106120 184600 106380
rect 184900 106120 185100 106380
rect 185400 106120 185600 106380
rect 185900 106120 186100 106380
rect 186400 106120 186600 106380
rect 186900 106120 187100 106380
rect 187400 106120 187600 106380
rect 187900 106120 188100 106380
rect 188400 106120 188600 106380
rect 188900 106120 189100 106380
rect 189400 106120 189600 106380
rect 189900 106120 190100 106380
rect 190400 106120 190600 106380
rect 190900 106120 191100 106380
rect 191400 106120 191600 106380
rect 191900 106120 192100 106380
rect 192400 106120 192600 106380
rect 192900 106120 193100 106380
rect 193400 106120 193600 106380
rect 193900 106120 194100 106380
rect 194400 106120 194600 106380
rect 194900 106120 195100 106380
rect 195400 106120 195600 106380
rect 195900 106120 196100 106380
rect 196400 106120 196600 106380
rect 196900 106120 197100 106380
rect 197400 106120 197600 106380
rect 197900 106120 198100 106380
rect 198400 106120 198600 106380
rect 198900 106120 199100 106380
rect 199400 106120 199600 106380
rect 199900 106120 200100 106380
rect 200400 106120 200600 106380
rect 200900 106120 201100 106380
rect 201400 106120 201600 106380
rect 201900 106120 202100 106380
rect 202400 106120 202600 106380
rect 202900 106120 203100 106380
rect 203400 106120 203600 106380
rect 203900 106120 204100 106380
rect 204400 106120 204600 106380
rect 204900 106120 205100 106380
rect 205400 106120 205600 106380
rect 205900 106120 206100 106380
rect 206400 106120 206600 106380
rect 206900 106120 207100 106380
rect 207400 106120 207600 106380
rect 207900 106120 208100 106380
rect 208400 106120 208600 106380
rect 208900 106120 209100 106380
rect 209400 106120 209600 106380
rect 209900 106120 210100 106380
rect 210400 106120 210600 106380
rect 210900 106120 211100 106380
rect 211400 106120 211600 106380
rect 211900 106120 212100 106380
rect 212400 106120 212600 106380
rect 212900 106120 213100 106380
rect 213400 106120 213600 106380
rect 213900 106120 214100 106380
rect 214400 106120 214600 106380
rect 214900 106120 215100 106380
rect 215400 106120 215600 106380
rect 215900 106120 216100 106380
rect 216400 106120 216600 106380
rect 216900 106120 217100 106380
rect 217400 106120 217600 106380
rect 217900 106120 218100 106380
rect 218400 106120 218600 106380
rect 218900 106120 219100 106380
rect 219400 106120 219600 106380
rect 219900 106120 220100 106380
rect 220400 106120 220600 106380
rect 220900 106120 221100 106380
rect 221400 106120 221600 106380
rect 221900 106120 222100 106380
rect 222400 106120 222600 106380
rect 222900 106120 223100 106380
rect 223400 106120 223600 106380
rect 223900 106120 224100 106380
rect 224400 106120 224600 106380
rect 224900 106120 225100 106380
rect 225400 106120 225600 106380
rect 225900 106120 226100 106380
rect 226400 106120 226600 106380
rect 226900 106120 227100 106380
rect 227400 106120 227600 106380
rect 227900 106120 228100 106380
rect 228400 106120 228600 106380
rect 228900 106120 229100 106380
rect 229400 106120 229600 106380
rect 229900 106120 230100 106380
rect 230400 106120 230600 106380
rect 230900 106120 231100 106380
rect 231400 106120 231600 106380
rect 231900 106120 232000 106380
rect 178000 106100 178120 106120
rect 178380 106100 178620 106120
rect 178880 106100 179120 106120
rect 179380 106100 179620 106120
rect 179880 106100 180120 106120
rect 180380 106100 180620 106120
rect 180880 106100 181120 106120
rect 181380 106100 181620 106120
rect 181880 106100 182120 106120
rect 182380 106100 182620 106120
rect 182880 106100 183120 106120
rect 183380 106100 183620 106120
rect 183880 106100 184120 106120
rect 184380 106100 184620 106120
rect 184880 106100 185120 106120
rect 185380 106100 185620 106120
rect 185880 106100 186120 106120
rect 186380 106100 186620 106120
rect 186880 106100 187120 106120
rect 187380 106100 187620 106120
rect 187880 106100 188120 106120
rect 188380 106100 188620 106120
rect 188880 106100 189120 106120
rect 189380 106100 189620 106120
rect 189880 106100 190120 106120
rect 190380 106100 190620 106120
rect 190880 106100 191120 106120
rect 191380 106100 191620 106120
rect 191880 106100 192120 106120
rect 192380 106100 192620 106120
rect 192880 106100 193120 106120
rect 193380 106100 193620 106120
rect 193880 106100 194120 106120
rect 194380 106100 194620 106120
rect 194880 106100 195120 106120
rect 195380 106100 195620 106120
rect 195880 106100 196120 106120
rect 196380 106100 196620 106120
rect 196880 106100 197120 106120
rect 197380 106100 197620 106120
rect 197880 106100 198120 106120
rect 198380 106100 198620 106120
rect 198880 106100 199120 106120
rect 199380 106100 199620 106120
rect 199880 106100 200120 106120
rect 200380 106100 200620 106120
rect 200880 106100 201120 106120
rect 201380 106100 201620 106120
rect 201880 106100 202120 106120
rect 202380 106100 202620 106120
rect 202880 106100 203120 106120
rect 203380 106100 203620 106120
rect 203880 106100 204120 106120
rect 204380 106100 204620 106120
rect 204880 106100 205120 106120
rect 205380 106100 205620 106120
rect 205880 106100 206120 106120
rect 206380 106100 206620 106120
rect 206880 106100 207120 106120
rect 207380 106100 207620 106120
rect 207880 106100 208120 106120
rect 208380 106100 208620 106120
rect 208880 106100 209120 106120
rect 209380 106100 209620 106120
rect 209880 106100 210120 106120
rect 210380 106100 210620 106120
rect 210880 106100 211120 106120
rect 211380 106100 211620 106120
rect 211880 106100 212120 106120
rect 212380 106100 212620 106120
rect 212880 106100 213120 106120
rect 213380 106100 213620 106120
rect 213880 106100 214120 106120
rect 214380 106100 214620 106120
rect 214880 106100 215120 106120
rect 215380 106100 215620 106120
rect 215880 106100 216120 106120
rect 216380 106100 216620 106120
rect 216880 106100 217120 106120
rect 217380 106100 217620 106120
rect 217880 106100 218120 106120
rect 218380 106100 218620 106120
rect 218880 106100 219120 106120
rect 219380 106100 219620 106120
rect 219880 106100 220120 106120
rect 220380 106100 220620 106120
rect 220880 106100 221120 106120
rect 221380 106100 221620 106120
rect 221880 106100 222120 106120
rect 222380 106100 222620 106120
rect 222880 106100 223120 106120
rect 223380 106100 223620 106120
rect 223880 106100 224120 106120
rect 224380 106100 224620 106120
rect 224880 106100 225120 106120
rect 225380 106100 225620 106120
rect 225880 106100 226120 106120
rect 226380 106100 226620 106120
rect 226880 106100 227120 106120
rect 227380 106100 227620 106120
rect 227880 106100 228120 106120
rect 228380 106100 228620 106120
rect 228880 106100 229120 106120
rect 229380 106100 229620 106120
rect 229880 106100 230120 106120
rect 230380 106100 230620 106120
rect 230880 106100 231120 106120
rect 231380 106100 231620 106120
rect 231880 106100 232000 106120
rect 178000 105900 232000 106100
rect 178000 105880 178120 105900
rect 178380 105880 178620 105900
rect 178880 105880 179120 105900
rect 179380 105880 179620 105900
rect 179880 105880 180120 105900
rect 180380 105880 180620 105900
rect 180880 105880 181120 105900
rect 181380 105880 181620 105900
rect 181880 105880 182120 105900
rect 182380 105880 182620 105900
rect 182880 105880 183120 105900
rect 183380 105880 183620 105900
rect 183880 105880 184120 105900
rect 184380 105880 184620 105900
rect 184880 105880 185120 105900
rect 185380 105880 185620 105900
rect 185880 105880 186120 105900
rect 186380 105880 186620 105900
rect 186880 105880 187120 105900
rect 187380 105880 187620 105900
rect 187880 105880 188120 105900
rect 188380 105880 188620 105900
rect 188880 105880 189120 105900
rect 189380 105880 189620 105900
rect 189880 105880 190120 105900
rect 190380 105880 190620 105900
rect 190880 105880 191120 105900
rect 191380 105880 191620 105900
rect 191880 105880 192120 105900
rect 192380 105880 192620 105900
rect 192880 105880 193120 105900
rect 193380 105880 193620 105900
rect 193880 105880 194120 105900
rect 194380 105880 194620 105900
rect 194880 105880 195120 105900
rect 195380 105880 195620 105900
rect 195880 105880 196120 105900
rect 196380 105880 196620 105900
rect 196880 105880 197120 105900
rect 197380 105880 197620 105900
rect 197880 105880 198120 105900
rect 198380 105880 198620 105900
rect 198880 105880 199120 105900
rect 199380 105880 199620 105900
rect 199880 105880 200120 105900
rect 200380 105880 200620 105900
rect 200880 105880 201120 105900
rect 201380 105880 201620 105900
rect 201880 105880 202120 105900
rect 202380 105880 202620 105900
rect 202880 105880 203120 105900
rect 203380 105880 203620 105900
rect 203880 105880 204120 105900
rect 204380 105880 204620 105900
rect 204880 105880 205120 105900
rect 205380 105880 205620 105900
rect 205880 105880 206120 105900
rect 206380 105880 206620 105900
rect 206880 105880 207120 105900
rect 207380 105880 207620 105900
rect 207880 105880 208120 105900
rect 208380 105880 208620 105900
rect 208880 105880 209120 105900
rect 209380 105880 209620 105900
rect 209880 105880 210120 105900
rect 210380 105880 210620 105900
rect 210880 105880 211120 105900
rect 211380 105880 211620 105900
rect 211880 105880 212120 105900
rect 212380 105880 212620 105900
rect 212880 105880 213120 105900
rect 213380 105880 213620 105900
rect 213880 105880 214120 105900
rect 214380 105880 214620 105900
rect 214880 105880 215120 105900
rect 215380 105880 215620 105900
rect 215880 105880 216120 105900
rect 216380 105880 216620 105900
rect 216880 105880 217120 105900
rect 217380 105880 217620 105900
rect 217880 105880 218120 105900
rect 218380 105880 218620 105900
rect 218880 105880 219120 105900
rect 219380 105880 219620 105900
rect 219880 105880 220120 105900
rect 220380 105880 220620 105900
rect 220880 105880 221120 105900
rect 221380 105880 221620 105900
rect 221880 105880 222120 105900
rect 222380 105880 222620 105900
rect 222880 105880 223120 105900
rect 223380 105880 223620 105900
rect 223880 105880 224120 105900
rect 224380 105880 224620 105900
rect 224880 105880 225120 105900
rect 225380 105880 225620 105900
rect 225880 105880 226120 105900
rect 226380 105880 226620 105900
rect 226880 105880 227120 105900
rect 227380 105880 227620 105900
rect 227880 105880 228120 105900
rect 228380 105880 228620 105900
rect 228880 105880 229120 105900
rect 229380 105880 229620 105900
rect 229880 105880 230120 105900
rect 230380 105880 230620 105900
rect 230880 105880 231120 105900
rect 231380 105880 231620 105900
rect 231880 105880 232000 105900
rect 178000 105620 178100 105880
rect 178400 105620 178600 105880
rect 178900 105620 179100 105880
rect 179400 105620 179600 105880
rect 179900 105620 180100 105880
rect 180400 105620 180600 105880
rect 180900 105620 181100 105880
rect 181400 105620 181600 105880
rect 181900 105620 182100 105880
rect 182400 105620 182600 105880
rect 182900 105620 183100 105880
rect 183400 105620 183600 105880
rect 183900 105620 184100 105880
rect 184400 105620 184600 105880
rect 184900 105620 185100 105880
rect 185400 105620 185600 105880
rect 185900 105620 186100 105880
rect 186400 105620 186600 105880
rect 186900 105620 187100 105880
rect 187400 105620 187600 105880
rect 187900 105620 188100 105880
rect 188400 105620 188600 105880
rect 188900 105620 189100 105880
rect 189400 105620 189600 105880
rect 189900 105620 190100 105880
rect 190400 105620 190600 105880
rect 190900 105620 191100 105880
rect 191400 105620 191600 105880
rect 191900 105620 192100 105880
rect 192400 105620 192600 105880
rect 192900 105620 193100 105880
rect 193400 105620 193600 105880
rect 193900 105620 194100 105880
rect 194400 105620 194600 105880
rect 194900 105620 195100 105880
rect 195400 105620 195600 105880
rect 195900 105620 196100 105880
rect 196400 105620 196600 105880
rect 196900 105620 197100 105880
rect 197400 105620 197600 105880
rect 197900 105620 198100 105880
rect 198400 105620 198600 105880
rect 198900 105620 199100 105880
rect 199400 105620 199600 105880
rect 199900 105620 200100 105880
rect 200400 105620 200600 105880
rect 200900 105620 201100 105880
rect 201400 105620 201600 105880
rect 201900 105620 202100 105880
rect 202400 105620 202600 105880
rect 202900 105620 203100 105880
rect 203400 105620 203600 105880
rect 203900 105620 204100 105880
rect 204400 105620 204600 105880
rect 204900 105620 205100 105880
rect 205400 105620 205600 105880
rect 205900 105620 206100 105880
rect 206400 105620 206600 105880
rect 206900 105620 207100 105880
rect 207400 105620 207600 105880
rect 207900 105620 208100 105880
rect 208400 105620 208600 105880
rect 208900 105620 209100 105880
rect 209400 105620 209600 105880
rect 209900 105620 210100 105880
rect 210400 105620 210600 105880
rect 210900 105620 211100 105880
rect 211400 105620 211600 105880
rect 211900 105620 212100 105880
rect 212400 105620 212600 105880
rect 212900 105620 213100 105880
rect 213400 105620 213600 105880
rect 213900 105620 214100 105880
rect 214400 105620 214600 105880
rect 214900 105620 215100 105880
rect 215400 105620 215600 105880
rect 215900 105620 216100 105880
rect 216400 105620 216600 105880
rect 216900 105620 217100 105880
rect 217400 105620 217600 105880
rect 217900 105620 218100 105880
rect 218400 105620 218600 105880
rect 218900 105620 219100 105880
rect 219400 105620 219600 105880
rect 219900 105620 220100 105880
rect 220400 105620 220600 105880
rect 220900 105620 221100 105880
rect 221400 105620 221600 105880
rect 221900 105620 222100 105880
rect 222400 105620 222600 105880
rect 222900 105620 223100 105880
rect 223400 105620 223600 105880
rect 223900 105620 224100 105880
rect 224400 105620 224600 105880
rect 224900 105620 225100 105880
rect 225400 105620 225600 105880
rect 225900 105620 226100 105880
rect 226400 105620 226600 105880
rect 226900 105620 227100 105880
rect 227400 105620 227600 105880
rect 227900 105620 228100 105880
rect 228400 105620 228600 105880
rect 228900 105620 229100 105880
rect 229400 105620 229600 105880
rect 229900 105620 230100 105880
rect 230400 105620 230600 105880
rect 230900 105620 231100 105880
rect 231400 105620 231600 105880
rect 231900 105620 232000 105880
rect 178000 105600 178120 105620
rect 178380 105600 178620 105620
rect 178880 105600 179120 105620
rect 179380 105600 179620 105620
rect 179880 105600 180120 105620
rect 180380 105600 180620 105620
rect 180880 105600 181120 105620
rect 181380 105600 181620 105620
rect 181880 105600 182120 105620
rect 182380 105600 182620 105620
rect 182880 105600 183120 105620
rect 183380 105600 183620 105620
rect 183880 105600 184120 105620
rect 184380 105600 184620 105620
rect 184880 105600 185120 105620
rect 185380 105600 185620 105620
rect 185880 105600 186120 105620
rect 186380 105600 186620 105620
rect 186880 105600 187120 105620
rect 187380 105600 187620 105620
rect 187880 105600 188120 105620
rect 188380 105600 188620 105620
rect 188880 105600 189120 105620
rect 189380 105600 189620 105620
rect 189880 105600 190120 105620
rect 190380 105600 190620 105620
rect 190880 105600 191120 105620
rect 191380 105600 191620 105620
rect 191880 105600 192120 105620
rect 192380 105600 192620 105620
rect 192880 105600 193120 105620
rect 193380 105600 193620 105620
rect 193880 105600 194120 105620
rect 194380 105600 194620 105620
rect 194880 105600 195120 105620
rect 195380 105600 195620 105620
rect 195880 105600 196120 105620
rect 196380 105600 196620 105620
rect 196880 105600 197120 105620
rect 197380 105600 197620 105620
rect 197880 105600 198120 105620
rect 198380 105600 198620 105620
rect 198880 105600 199120 105620
rect 199380 105600 199620 105620
rect 199880 105600 200120 105620
rect 200380 105600 200620 105620
rect 200880 105600 201120 105620
rect 201380 105600 201620 105620
rect 201880 105600 202120 105620
rect 202380 105600 202620 105620
rect 202880 105600 203120 105620
rect 203380 105600 203620 105620
rect 203880 105600 204120 105620
rect 204380 105600 204620 105620
rect 204880 105600 205120 105620
rect 205380 105600 205620 105620
rect 205880 105600 206120 105620
rect 206380 105600 206620 105620
rect 206880 105600 207120 105620
rect 207380 105600 207620 105620
rect 207880 105600 208120 105620
rect 208380 105600 208620 105620
rect 208880 105600 209120 105620
rect 209380 105600 209620 105620
rect 209880 105600 210120 105620
rect 210380 105600 210620 105620
rect 210880 105600 211120 105620
rect 211380 105600 211620 105620
rect 211880 105600 212120 105620
rect 212380 105600 212620 105620
rect 212880 105600 213120 105620
rect 213380 105600 213620 105620
rect 213880 105600 214120 105620
rect 214380 105600 214620 105620
rect 214880 105600 215120 105620
rect 215380 105600 215620 105620
rect 215880 105600 216120 105620
rect 216380 105600 216620 105620
rect 216880 105600 217120 105620
rect 217380 105600 217620 105620
rect 217880 105600 218120 105620
rect 218380 105600 218620 105620
rect 218880 105600 219120 105620
rect 219380 105600 219620 105620
rect 219880 105600 220120 105620
rect 220380 105600 220620 105620
rect 220880 105600 221120 105620
rect 221380 105600 221620 105620
rect 221880 105600 222120 105620
rect 222380 105600 222620 105620
rect 222880 105600 223120 105620
rect 223380 105600 223620 105620
rect 223880 105600 224120 105620
rect 224380 105600 224620 105620
rect 224880 105600 225120 105620
rect 225380 105600 225620 105620
rect 225880 105600 226120 105620
rect 226380 105600 226620 105620
rect 226880 105600 227120 105620
rect 227380 105600 227620 105620
rect 227880 105600 228120 105620
rect 228380 105600 228620 105620
rect 228880 105600 229120 105620
rect 229380 105600 229620 105620
rect 229880 105600 230120 105620
rect 230380 105600 230620 105620
rect 230880 105600 231120 105620
rect 231380 105600 231620 105620
rect 231880 105600 232000 105620
rect 178000 105400 232000 105600
rect 178000 105380 178120 105400
rect 178380 105380 178620 105400
rect 178880 105380 179120 105400
rect 179380 105380 179620 105400
rect 179880 105380 180120 105400
rect 180380 105380 180620 105400
rect 180880 105380 181120 105400
rect 181380 105380 181620 105400
rect 181880 105380 182120 105400
rect 182380 105380 182620 105400
rect 182880 105380 183120 105400
rect 183380 105380 183620 105400
rect 183880 105380 184120 105400
rect 184380 105380 184620 105400
rect 184880 105380 185120 105400
rect 185380 105380 185620 105400
rect 185880 105380 186120 105400
rect 186380 105380 186620 105400
rect 186880 105380 187120 105400
rect 187380 105380 187620 105400
rect 187880 105380 188120 105400
rect 188380 105380 188620 105400
rect 188880 105380 189120 105400
rect 189380 105380 189620 105400
rect 189880 105380 190120 105400
rect 190380 105380 190620 105400
rect 190880 105380 191120 105400
rect 191380 105380 191620 105400
rect 191880 105380 192120 105400
rect 192380 105380 192620 105400
rect 192880 105380 193120 105400
rect 193380 105380 193620 105400
rect 193880 105380 194120 105400
rect 194380 105380 194620 105400
rect 194880 105380 195120 105400
rect 195380 105380 195620 105400
rect 195880 105380 196120 105400
rect 196380 105380 196620 105400
rect 196880 105380 197120 105400
rect 197380 105380 197620 105400
rect 197880 105380 198120 105400
rect 198380 105380 198620 105400
rect 198880 105380 199120 105400
rect 199380 105380 199620 105400
rect 199880 105380 200120 105400
rect 200380 105380 200620 105400
rect 200880 105380 201120 105400
rect 201380 105380 201620 105400
rect 201880 105380 202120 105400
rect 202380 105380 202620 105400
rect 202880 105380 203120 105400
rect 203380 105380 203620 105400
rect 203880 105380 204120 105400
rect 204380 105380 204620 105400
rect 204880 105380 205120 105400
rect 205380 105380 205620 105400
rect 205880 105380 206120 105400
rect 206380 105380 206620 105400
rect 206880 105380 207120 105400
rect 207380 105380 207620 105400
rect 207880 105380 208120 105400
rect 208380 105380 208620 105400
rect 208880 105380 209120 105400
rect 209380 105380 209620 105400
rect 209880 105380 210120 105400
rect 210380 105380 210620 105400
rect 210880 105380 211120 105400
rect 211380 105380 211620 105400
rect 211880 105380 212120 105400
rect 212380 105380 212620 105400
rect 212880 105380 213120 105400
rect 213380 105380 213620 105400
rect 213880 105380 214120 105400
rect 214380 105380 214620 105400
rect 214880 105380 215120 105400
rect 215380 105380 215620 105400
rect 215880 105380 216120 105400
rect 216380 105380 216620 105400
rect 216880 105380 217120 105400
rect 217380 105380 217620 105400
rect 217880 105380 218120 105400
rect 218380 105380 218620 105400
rect 218880 105380 219120 105400
rect 219380 105380 219620 105400
rect 219880 105380 220120 105400
rect 220380 105380 220620 105400
rect 220880 105380 221120 105400
rect 221380 105380 221620 105400
rect 221880 105380 222120 105400
rect 222380 105380 222620 105400
rect 222880 105380 223120 105400
rect 223380 105380 223620 105400
rect 223880 105380 224120 105400
rect 224380 105380 224620 105400
rect 224880 105380 225120 105400
rect 225380 105380 225620 105400
rect 225880 105380 226120 105400
rect 226380 105380 226620 105400
rect 226880 105380 227120 105400
rect 227380 105380 227620 105400
rect 227880 105380 228120 105400
rect 228380 105380 228620 105400
rect 228880 105380 229120 105400
rect 229380 105380 229620 105400
rect 229880 105380 230120 105400
rect 230380 105380 230620 105400
rect 230880 105380 231120 105400
rect 231380 105380 231620 105400
rect 231880 105380 232000 105400
rect 178000 105120 178100 105380
rect 178400 105120 178600 105380
rect 178900 105120 179100 105380
rect 179400 105120 179600 105380
rect 179900 105120 180100 105380
rect 180400 105120 180600 105380
rect 180900 105120 181100 105380
rect 181400 105120 181600 105380
rect 181900 105120 182100 105380
rect 182400 105120 182600 105380
rect 182900 105120 183100 105380
rect 183400 105120 183600 105380
rect 183900 105120 184100 105380
rect 184400 105120 184600 105380
rect 184900 105120 185100 105380
rect 185400 105120 185600 105380
rect 185900 105120 186100 105380
rect 186400 105120 186600 105380
rect 186900 105120 187100 105380
rect 187400 105120 187600 105380
rect 187900 105120 188100 105380
rect 188400 105120 188600 105380
rect 188900 105120 189100 105380
rect 189400 105120 189600 105380
rect 189900 105120 190100 105380
rect 190400 105120 190600 105380
rect 190900 105120 191100 105380
rect 191400 105120 191600 105380
rect 191900 105120 192100 105380
rect 192400 105120 192600 105380
rect 192900 105120 193100 105380
rect 193400 105120 193600 105380
rect 193900 105120 194100 105380
rect 194400 105120 194600 105380
rect 194900 105120 195100 105380
rect 195400 105120 195600 105380
rect 195900 105120 196100 105380
rect 196400 105120 196600 105380
rect 196900 105120 197100 105380
rect 197400 105120 197600 105380
rect 197900 105120 198100 105380
rect 198400 105120 198600 105380
rect 198900 105120 199100 105380
rect 199400 105120 199600 105380
rect 199900 105120 200100 105380
rect 200400 105120 200600 105380
rect 200900 105120 201100 105380
rect 201400 105120 201600 105380
rect 201900 105120 202100 105380
rect 202400 105120 202600 105380
rect 202900 105120 203100 105380
rect 203400 105120 203600 105380
rect 203900 105120 204100 105380
rect 204400 105120 204600 105380
rect 204900 105120 205100 105380
rect 205400 105120 205600 105380
rect 205900 105120 206100 105380
rect 206400 105120 206600 105380
rect 206900 105120 207100 105380
rect 207400 105120 207600 105380
rect 207900 105120 208100 105380
rect 208400 105120 208600 105380
rect 208900 105120 209100 105380
rect 209400 105120 209600 105380
rect 209900 105120 210100 105380
rect 210400 105120 210600 105380
rect 210900 105120 211100 105380
rect 211400 105120 211600 105380
rect 211900 105120 212100 105380
rect 212400 105120 212600 105380
rect 212900 105120 213100 105380
rect 213400 105120 213600 105380
rect 213900 105120 214100 105380
rect 214400 105120 214600 105380
rect 214900 105120 215100 105380
rect 215400 105120 215600 105380
rect 215900 105120 216100 105380
rect 216400 105120 216600 105380
rect 216900 105120 217100 105380
rect 217400 105120 217600 105380
rect 217900 105120 218100 105380
rect 218400 105120 218600 105380
rect 218900 105120 219100 105380
rect 219400 105120 219600 105380
rect 219900 105120 220100 105380
rect 220400 105120 220600 105380
rect 220900 105120 221100 105380
rect 221400 105120 221600 105380
rect 221900 105120 222100 105380
rect 222400 105120 222600 105380
rect 222900 105120 223100 105380
rect 223400 105120 223600 105380
rect 223900 105120 224100 105380
rect 224400 105120 224600 105380
rect 224900 105120 225100 105380
rect 225400 105120 225600 105380
rect 225900 105120 226100 105380
rect 226400 105120 226600 105380
rect 226900 105120 227100 105380
rect 227400 105120 227600 105380
rect 227900 105120 228100 105380
rect 228400 105120 228600 105380
rect 228900 105120 229100 105380
rect 229400 105120 229600 105380
rect 229900 105120 230100 105380
rect 230400 105120 230600 105380
rect 230900 105120 231100 105380
rect 231400 105120 231600 105380
rect 231900 105120 232000 105380
rect 178000 105100 178120 105120
rect 178380 105100 178620 105120
rect 178880 105100 179120 105120
rect 179380 105100 179620 105120
rect 179880 105100 180120 105120
rect 180380 105100 180620 105120
rect 180880 105100 181120 105120
rect 181380 105100 181620 105120
rect 181880 105100 182120 105120
rect 182380 105100 182620 105120
rect 182880 105100 183120 105120
rect 183380 105100 183620 105120
rect 183880 105100 184120 105120
rect 184380 105100 184620 105120
rect 184880 105100 185120 105120
rect 185380 105100 185620 105120
rect 185880 105100 186120 105120
rect 186380 105100 186620 105120
rect 186880 105100 187120 105120
rect 187380 105100 187620 105120
rect 187880 105100 188120 105120
rect 188380 105100 188620 105120
rect 188880 105100 189120 105120
rect 189380 105100 189620 105120
rect 189880 105100 190120 105120
rect 190380 105100 190620 105120
rect 190880 105100 191120 105120
rect 191380 105100 191620 105120
rect 191880 105100 192120 105120
rect 192380 105100 192620 105120
rect 192880 105100 193120 105120
rect 193380 105100 193620 105120
rect 193880 105100 194120 105120
rect 194380 105100 194620 105120
rect 194880 105100 195120 105120
rect 195380 105100 195620 105120
rect 195880 105100 196120 105120
rect 196380 105100 196620 105120
rect 196880 105100 197120 105120
rect 197380 105100 197620 105120
rect 197880 105100 198120 105120
rect 198380 105100 198620 105120
rect 198880 105100 199120 105120
rect 199380 105100 199620 105120
rect 199880 105100 200120 105120
rect 200380 105100 200620 105120
rect 200880 105100 201120 105120
rect 201380 105100 201620 105120
rect 201880 105100 202120 105120
rect 202380 105100 202620 105120
rect 202880 105100 203120 105120
rect 203380 105100 203620 105120
rect 203880 105100 204120 105120
rect 204380 105100 204620 105120
rect 204880 105100 205120 105120
rect 205380 105100 205620 105120
rect 205880 105100 206120 105120
rect 206380 105100 206620 105120
rect 206880 105100 207120 105120
rect 207380 105100 207620 105120
rect 207880 105100 208120 105120
rect 208380 105100 208620 105120
rect 208880 105100 209120 105120
rect 209380 105100 209620 105120
rect 209880 105100 210120 105120
rect 210380 105100 210620 105120
rect 210880 105100 211120 105120
rect 211380 105100 211620 105120
rect 211880 105100 212120 105120
rect 212380 105100 212620 105120
rect 212880 105100 213120 105120
rect 213380 105100 213620 105120
rect 213880 105100 214120 105120
rect 214380 105100 214620 105120
rect 214880 105100 215120 105120
rect 215380 105100 215620 105120
rect 215880 105100 216120 105120
rect 216380 105100 216620 105120
rect 216880 105100 217120 105120
rect 217380 105100 217620 105120
rect 217880 105100 218120 105120
rect 218380 105100 218620 105120
rect 218880 105100 219120 105120
rect 219380 105100 219620 105120
rect 219880 105100 220120 105120
rect 220380 105100 220620 105120
rect 220880 105100 221120 105120
rect 221380 105100 221620 105120
rect 221880 105100 222120 105120
rect 222380 105100 222620 105120
rect 222880 105100 223120 105120
rect 223380 105100 223620 105120
rect 223880 105100 224120 105120
rect 224380 105100 224620 105120
rect 224880 105100 225120 105120
rect 225380 105100 225620 105120
rect 225880 105100 226120 105120
rect 226380 105100 226620 105120
rect 226880 105100 227120 105120
rect 227380 105100 227620 105120
rect 227880 105100 228120 105120
rect 228380 105100 228620 105120
rect 228880 105100 229120 105120
rect 229380 105100 229620 105120
rect 229880 105100 230120 105120
rect 230380 105100 230620 105120
rect 230880 105100 231120 105120
rect 231380 105100 231620 105120
rect 231880 105100 232000 105120
rect 178000 104900 232000 105100
rect 178000 104880 178120 104900
rect 178380 104880 178620 104900
rect 178880 104880 179120 104900
rect 179380 104880 179620 104900
rect 179880 104880 180120 104900
rect 180380 104880 180620 104900
rect 180880 104880 181120 104900
rect 181380 104880 181620 104900
rect 181880 104880 182120 104900
rect 182380 104880 182620 104900
rect 182880 104880 183120 104900
rect 183380 104880 183620 104900
rect 183880 104880 184120 104900
rect 184380 104880 184620 104900
rect 184880 104880 185120 104900
rect 185380 104880 185620 104900
rect 185880 104880 186120 104900
rect 186380 104880 186620 104900
rect 186880 104880 187120 104900
rect 187380 104880 187620 104900
rect 187880 104880 188120 104900
rect 188380 104880 188620 104900
rect 188880 104880 189120 104900
rect 189380 104880 189620 104900
rect 189880 104880 190120 104900
rect 190380 104880 190620 104900
rect 190880 104880 191120 104900
rect 191380 104880 191620 104900
rect 191880 104880 192120 104900
rect 192380 104880 192620 104900
rect 192880 104880 193120 104900
rect 193380 104880 193620 104900
rect 193880 104880 194120 104900
rect 194380 104880 194620 104900
rect 194880 104880 195120 104900
rect 195380 104880 195620 104900
rect 195880 104880 196120 104900
rect 196380 104880 196620 104900
rect 196880 104880 197120 104900
rect 197380 104880 197620 104900
rect 197880 104880 198120 104900
rect 198380 104880 198620 104900
rect 198880 104880 199120 104900
rect 199380 104880 199620 104900
rect 199880 104880 200120 104900
rect 200380 104880 200620 104900
rect 200880 104880 201120 104900
rect 201380 104880 201620 104900
rect 201880 104880 202120 104900
rect 202380 104880 202620 104900
rect 202880 104880 203120 104900
rect 203380 104880 203620 104900
rect 203880 104880 204120 104900
rect 204380 104880 204620 104900
rect 204880 104880 205120 104900
rect 205380 104880 205620 104900
rect 205880 104880 206120 104900
rect 206380 104880 206620 104900
rect 206880 104880 207120 104900
rect 207380 104880 207620 104900
rect 207880 104880 208120 104900
rect 208380 104880 208620 104900
rect 208880 104880 209120 104900
rect 209380 104880 209620 104900
rect 209880 104880 210120 104900
rect 210380 104880 210620 104900
rect 210880 104880 211120 104900
rect 211380 104880 211620 104900
rect 211880 104880 212120 104900
rect 212380 104880 212620 104900
rect 212880 104880 213120 104900
rect 213380 104880 213620 104900
rect 213880 104880 214120 104900
rect 214380 104880 214620 104900
rect 214880 104880 215120 104900
rect 215380 104880 215620 104900
rect 215880 104880 216120 104900
rect 216380 104880 216620 104900
rect 216880 104880 217120 104900
rect 217380 104880 217620 104900
rect 217880 104880 218120 104900
rect 218380 104880 218620 104900
rect 218880 104880 219120 104900
rect 219380 104880 219620 104900
rect 219880 104880 220120 104900
rect 220380 104880 220620 104900
rect 220880 104880 221120 104900
rect 221380 104880 221620 104900
rect 221880 104880 222120 104900
rect 222380 104880 222620 104900
rect 222880 104880 223120 104900
rect 223380 104880 223620 104900
rect 223880 104880 224120 104900
rect 224380 104880 224620 104900
rect 224880 104880 225120 104900
rect 225380 104880 225620 104900
rect 225880 104880 226120 104900
rect 226380 104880 226620 104900
rect 226880 104880 227120 104900
rect 227380 104880 227620 104900
rect 227880 104880 228120 104900
rect 228380 104880 228620 104900
rect 228880 104880 229120 104900
rect 229380 104880 229620 104900
rect 229880 104880 230120 104900
rect 230380 104880 230620 104900
rect 230880 104880 231120 104900
rect 231380 104880 231620 104900
rect 231880 104880 232000 104900
rect 178000 104620 178100 104880
rect 178400 104620 178600 104880
rect 178900 104620 179100 104880
rect 179400 104620 179600 104880
rect 179900 104620 180100 104880
rect 180400 104620 180600 104880
rect 180900 104620 181100 104880
rect 181400 104620 181600 104880
rect 181900 104620 182100 104880
rect 182400 104620 182600 104880
rect 182900 104620 183100 104880
rect 183400 104620 183600 104880
rect 183900 104620 184100 104880
rect 184400 104620 184600 104880
rect 184900 104620 185100 104880
rect 185400 104620 185600 104880
rect 185900 104620 186100 104880
rect 186400 104620 186600 104880
rect 186900 104620 187100 104880
rect 187400 104620 187600 104880
rect 187900 104620 188100 104880
rect 188400 104620 188600 104880
rect 188900 104620 189100 104880
rect 189400 104620 189600 104880
rect 189900 104620 190100 104880
rect 190400 104620 190600 104880
rect 190900 104620 191100 104880
rect 191400 104620 191600 104880
rect 191900 104620 192100 104880
rect 192400 104620 192600 104880
rect 192900 104620 193100 104880
rect 193400 104620 193600 104880
rect 193900 104620 194100 104880
rect 194400 104620 194600 104880
rect 194900 104620 195100 104880
rect 195400 104620 195600 104880
rect 195900 104620 196100 104880
rect 196400 104620 196600 104880
rect 196900 104620 197100 104880
rect 197400 104620 197600 104880
rect 197900 104620 198100 104880
rect 198400 104620 198600 104880
rect 198900 104620 199100 104880
rect 199400 104620 199600 104880
rect 199900 104620 200100 104880
rect 200400 104620 200600 104880
rect 200900 104620 201100 104880
rect 201400 104620 201600 104880
rect 201900 104620 202100 104880
rect 202400 104620 202600 104880
rect 202900 104620 203100 104880
rect 203400 104620 203600 104880
rect 203900 104620 204100 104880
rect 204400 104620 204600 104880
rect 204900 104620 205100 104880
rect 205400 104620 205600 104880
rect 205900 104620 206100 104880
rect 206400 104620 206600 104880
rect 206900 104620 207100 104880
rect 207400 104620 207600 104880
rect 207900 104620 208100 104880
rect 208400 104620 208600 104880
rect 208900 104620 209100 104880
rect 209400 104620 209600 104880
rect 209900 104620 210100 104880
rect 210400 104620 210600 104880
rect 210900 104620 211100 104880
rect 211400 104620 211600 104880
rect 211900 104620 212100 104880
rect 212400 104620 212600 104880
rect 212900 104620 213100 104880
rect 213400 104620 213600 104880
rect 213900 104620 214100 104880
rect 214400 104620 214600 104880
rect 214900 104620 215100 104880
rect 215400 104620 215600 104880
rect 215900 104620 216100 104880
rect 216400 104620 216600 104880
rect 216900 104620 217100 104880
rect 217400 104620 217600 104880
rect 217900 104620 218100 104880
rect 218400 104620 218600 104880
rect 218900 104620 219100 104880
rect 219400 104620 219600 104880
rect 219900 104620 220100 104880
rect 220400 104620 220600 104880
rect 220900 104620 221100 104880
rect 221400 104620 221600 104880
rect 221900 104620 222100 104880
rect 222400 104620 222600 104880
rect 222900 104620 223100 104880
rect 223400 104620 223600 104880
rect 223900 104620 224100 104880
rect 224400 104620 224600 104880
rect 224900 104620 225100 104880
rect 225400 104620 225600 104880
rect 225900 104620 226100 104880
rect 226400 104620 226600 104880
rect 226900 104620 227100 104880
rect 227400 104620 227600 104880
rect 227900 104620 228100 104880
rect 228400 104620 228600 104880
rect 228900 104620 229100 104880
rect 229400 104620 229600 104880
rect 229900 104620 230100 104880
rect 230400 104620 230600 104880
rect 230900 104620 231100 104880
rect 231400 104620 231600 104880
rect 231900 104620 232000 104880
rect 178000 104600 178120 104620
rect 178380 104600 178620 104620
rect 178880 104600 179120 104620
rect 179380 104600 179620 104620
rect 179880 104600 180120 104620
rect 180380 104600 180620 104620
rect 180880 104600 181120 104620
rect 181380 104600 181620 104620
rect 181880 104600 182120 104620
rect 182380 104600 182620 104620
rect 182880 104600 183120 104620
rect 183380 104600 183620 104620
rect 183880 104600 184120 104620
rect 184380 104600 184620 104620
rect 184880 104600 185120 104620
rect 185380 104600 185620 104620
rect 185880 104600 186120 104620
rect 186380 104600 186620 104620
rect 186880 104600 187120 104620
rect 187380 104600 187620 104620
rect 187880 104600 188120 104620
rect 188380 104600 188620 104620
rect 188880 104600 189120 104620
rect 189380 104600 189620 104620
rect 189880 104600 190120 104620
rect 190380 104600 190620 104620
rect 190880 104600 191120 104620
rect 191380 104600 191620 104620
rect 191880 104600 192120 104620
rect 192380 104600 192620 104620
rect 192880 104600 193120 104620
rect 193380 104600 193620 104620
rect 193880 104600 194120 104620
rect 194380 104600 194620 104620
rect 194880 104600 195120 104620
rect 195380 104600 195620 104620
rect 195880 104600 196120 104620
rect 196380 104600 196620 104620
rect 196880 104600 197120 104620
rect 197380 104600 197620 104620
rect 197880 104600 198120 104620
rect 198380 104600 198620 104620
rect 198880 104600 199120 104620
rect 199380 104600 199620 104620
rect 199880 104600 200120 104620
rect 200380 104600 200620 104620
rect 200880 104600 201120 104620
rect 201380 104600 201620 104620
rect 201880 104600 202120 104620
rect 202380 104600 202620 104620
rect 202880 104600 203120 104620
rect 203380 104600 203620 104620
rect 203880 104600 204120 104620
rect 204380 104600 204620 104620
rect 204880 104600 205120 104620
rect 205380 104600 205620 104620
rect 205880 104600 206120 104620
rect 206380 104600 206620 104620
rect 206880 104600 207120 104620
rect 207380 104600 207620 104620
rect 207880 104600 208120 104620
rect 208380 104600 208620 104620
rect 208880 104600 209120 104620
rect 209380 104600 209620 104620
rect 209880 104600 210120 104620
rect 210380 104600 210620 104620
rect 210880 104600 211120 104620
rect 211380 104600 211620 104620
rect 211880 104600 212120 104620
rect 212380 104600 212620 104620
rect 212880 104600 213120 104620
rect 213380 104600 213620 104620
rect 213880 104600 214120 104620
rect 214380 104600 214620 104620
rect 214880 104600 215120 104620
rect 215380 104600 215620 104620
rect 215880 104600 216120 104620
rect 216380 104600 216620 104620
rect 216880 104600 217120 104620
rect 217380 104600 217620 104620
rect 217880 104600 218120 104620
rect 218380 104600 218620 104620
rect 218880 104600 219120 104620
rect 219380 104600 219620 104620
rect 219880 104600 220120 104620
rect 220380 104600 220620 104620
rect 220880 104600 221120 104620
rect 221380 104600 221620 104620
rect 221880 104600 222120 104620
rect 222380 104600 222620 104620
rect 222880 104600 223120 104620
rect 223380 104600 223620 104620
rect 223880 104600 224120 104620
rect 224380 104600 224620 104620
rect 224880 104600 225120 104620
rect 225380 104600 225620 104620
rect 225880 104600 226120 104620
rect 226380 104600 226620 104620
rect 226880 104600 227120 104620
rect 227380 104600 227620 104620
rect 227880 104600 228120 104620
rect 228380 104600 228620 104620
rect 228880 104600 229120 104620
rect 229380 104600 229620 104620
rect 229880 104600 230120 104620
rect 230380 104600 230620 104620
rect 230880 104600 231120 104620
rect 231380 104600 231620 104620
rect 231880 104600 232000 104620
rect 178000 104400 232000 104600
rect 178000 104380 178120 104400
rect 178380 104380 178620 104400
rect 178880 104380 179120 104400
rect 179380 104380 179620 104400
rect 179880 104380 180120 104400
rect 180380 104380 180620 104400
rect 180880 104380 181120 104400
rect 181380 104380 181620 104400
rect 181880 104380 182120 104400
rect 182380 104380 182620 104400
rect 182880 104380 183120 104400
rect 183380 104380 183620 104400
rect 183880 104380 184120 104400
rect 184380 104380 184620 104400
rect 184880 104380 185120 104400
rect 185380 104380 185620 104400
rect 185880 104380 186120 104400
rect 186380 104380 186620 104400
rect 186880 104380 187120 104400
rect 187380 104380 187620 104400
rect 187880 104380 188120 104400
rect 188380 104380 188620 104400
rect 188880 104380 189120 104400
rect 189380 104380 189620 104400
rect 189880 104380 190120 104400
rect 190380 104380 190620 104400
rect 190880 104380 191120 104400
rect 191380 104380 191620 104400
rect 191880 104380 192120 104400
rect 192380 104380 192620 104400
rect 192880 104380 193120 104400
rect 193380 104380 193620 104400
rect 193880 104380 194120 104400
rect 194380 104380 194620 104400
rect 194880 104380 195120 104400
rect 195380 104380 195620 104400
rect 195880 104380 196120 104400
rect 196380 104380 196620 104400
rect 196880 104380 197120 104400
rect 197380 104380 197620 104400
rect 197880 104380 198120 104400
rect 198380 104380 198620 104400
rect 198880 104380 199120 104400
rect 199380 104380 199620 104400
rect 199880 104380 200120 104400
rect 200380 104380 200620 104400
rect 200880 104380 201120 104400
rect 201380 104380 201620 104400
rect 201880 104380 202120 104400
rect 202380 104380 202620 104400
rect 202880 104380 203120 104400
rect 203380 104380 203620 104400
rect 203880 104380 204120 104400
rect 204380 104380 204620 104400
rect 204880 104380 205120 104400
rect 205380 104380 205620 104400
rect 205880 104380 206120 104400
rect 206380 104380 206620 104400
rect 206880 104380 207120 104400
rect 207380 104380 207620 104400
rect 207880 104380 208120 104400
rect 208380 104380 208620 104400
rect 208880 104380 209120 104400
rect 209380 104380 209620 104400
rect 209880 104380 210120 104400
rect 210380 104380 210620 104400
rect 210880 104380 211120 104400
rect 211380 104380 211620 104400
rect 211880 104380 212120 104400
rect 212380 104380 212620 104400
rect 212880 104380 213120 104400
rect 213380 104380 213620 104400
rect 213880 104380 214120 104400
rect 214380 104380 214620 104400
rect 214880 104380 215120 104400
rect 215380 104380 215620 104400
rect 215880 104380 216120 104400
rect 216380 104380 216620 104400
rect 216880 104380 217120 104400
rect 217380 104380 217620 104400
rect 217880 104380 218120 104400
rect 218380 104380 218620 104400
rect 218880 104380 219120 104400
rect 219380 104380 219620 104400
rect 219880 104380 220120 104400
rect 220380 104380 220620 104400
rect 220880 104380 221120 104400
rect 221380 104380 221620 104400
rect 221880 104380 222120 104400
rect 222380 104380 222620 104400
rect 222880 104380 223120 104400
rect 223380 104380 223620 104400
rect 223880 104380 224120 104400
rect 224380 104380 224620 104400
rect 224880 104380 225120 104400
rect 225380 104380 225620 104400
rect 225880 104380 226120 104400
rect 226380 104380 226620 104400
rect 226880 104380 227120 104400
rect 227380 104380 227620 104400
rect 227880 104380 228120 104400
rect 228380 104380 228620 104400
rect 228880 104380 229120 104400
rect 229380 104380 229620 104400
rect 229880 104380 230120 104400
rect 230380 104380 230620 104400
rect 230880 104380 231120 104400
rect 231380 104380 231620 104400
rect 231880 104380 232000 104400
rect 178000 104120 178100 104380
rect 178400 104120 178600 104380
rect 178900 104120 179100 104380
rect 179400 104120 179600 104380
rect 179900 104120 180100 104380
rect 180400 104120 180600 104380
rect 180900 104120 181100 104380
rect 181400 104120 181600 104380
rect 181900 104120 182100 104380
rect 182400 104120 182600 104380
rect 182900 104120 183100 104380
rect 183400 104120 183600 104380
rect 183900 104120 184100 104380
rect 184400 104120 184600 104380
rect 184900 104120 185100 104380
rect 185400 104120 185600 104380
rect 185900 104120 186100 104380
rect 186400 104120 186600 104380
rect 186900 104120 187100 104380
rect 187400 104120 187600 104380
rect 187900 104120 188100 104380
rect 188400 104120 188600 104380
rect 188900 104120 189100 104380
rect 189400 104120 189600 104380
rect 189900 104120 190100 104380
rect 190400 104120 190600 104380
rect 190900 104120 191100 104380
rect 191400 104120 191600 104380
rect 191900 104120 192100 104380
rect 192400 104120 192600 104380
rect 192900 104120 193100 104380
rect 193400 104120 193600 104380
rect 193900 104120 194100 104380
rect 194400 104120 194600 104380
rect 194900 104120 195100 104380
rect 195400 104120 195600 104380
rect 195900 104120 196100 104380
rect 196400 104120 196600 104380
rect 196900 104120 197100 104380
rect 197400 104120 197600 104380
rect 197900 104120 198100 104380
rect 198400 104120 198600 104380
rect 198900 104120 199100 104380
rect 199400 104120 199600 104380
rect 199900 104120 200100 104380
rect 200400 104120 200600 104380
rect 200900 104120 201100 104380
rect 201400 104120 201600 104380
rect 201900 104120 202100 104380
rect 202400 104120 202600 104380
rect 202900 104120 203100 104380
rect 203400 104120 203600 104380
rect 203900 104120 204100 104380
rect 204400 104120 204600 104380
rect 204900 104120 205100 104380
rect 205400 104120 205600 104380
rect 205900 104120 206100 104380
rect 206400 104120 206600 104380
rect 206900 104120 207100 104380
rect 207400 104120 207600 104380
rect 207900 104120 208100 104380
rect 208400 104120 208600 104380
rect 208900 104120 209100 104380
rect 209400 104120 209600 104380
rect 209900 104120 210100 104380
rect 210400 104120 210600 104380
rect 210900 104120 211100 104380
rect 211400 104120 211600 104380
rect 211900 104120 212100 104380
rect 212400 104120 212600 104380
rect 212900 104120 213100 104380
rect 213400 104120 213600 104380
rect 213900 104120 214100 104380
rect 214400 104120 214600 104380
rect 214900 104120 215100 104380
rect 215400 104120 215600 104380
rect 215900 104120 216100 104380
rect 216400 104120 216600 104380
rect 216900 104120 217100 104380
rect 217400 104120 217600 104380
rect 217900 104120 218100 104380
rect 218400 104120 218600 104380
rect 218900 104120 219100 104380
rect 219400 104120 219600 104380
rect 219900 104120 220100 104380
rect 220400 104120 220600 104380
rect 220900 104120 221100 104380
rect 221400 104120 221600 104380
rect 221900 104120 222100 104380
rect 222400 104120 222600 104380
rect 222900 104120 223100 104380
rect 223400 104120 223600 104380
rect 223900 104120 224100 104380
rect 224400 104120 224600 104380
rect 224900 104120 225100 104380
rect 225400 104120 225600 104380
rect 225900 104120 226100 104380
rect 226400 104120 226600 104380
rect 226900 104120 227100 104380
rect 227400 104120 227600 104380
rect 227900 104120 228100 104380
rect 228400 104120 228600 104380
rect 228900 104120 229100 104380
rect 229400 104120 229600 104380
rect 229900 104120 230100 104380
rect 230400 104120 230600 104380
rect 230900 104120 231100 104380
rect 231400 104120 231600 104380
rect 231900 104120 232000 104380
rect 178000 104100 178120 104120
rect 178380 104100 178620 104120
rect 178880 104100 179120 104120
rect 179380 104100 179620 104120
rect 179880 104100 180120 104120
rect 180380 104100 180620 104120
rect 180880 104100 181120 104120
rect 181380 104100 181620 104120
rect 181880 104100 182120 104120
rect 182380 104100 182620 104120
rect 182880 104100 183120 104120
rect 183380 104100 183620 104120
rect 183880 104100 184120 104120
rect 184380 104100 184620 104120
rect 184880 104100 185120 104120
rect 185380 104100 185620 104120
rect 185880 104100 186120 104120
rect 186380 104100 186620 104120
rect 186880 104100 187120 104120
rect 187380 104100 187620 104120
rect 187880 104100 188120 104120
rect 188380 104100 188620 104120
rect 188880 104100 189120 104120
rect 189380 104100 189620 104120
rect 189880 104100 190120 104120
rect 190380 104100 190620 104120
rect 190880 104100 191120 104120
rect 191380 104100 191620 104120
rect 191880 104100 192120 104120
rect 192380 104100 192620 104120
rect 192880 104100 193120 104120
rect 193380 104100 193620 104120
rect 193880 104100 194120 104120
rect 194380 104100 194620 104120
rect 194880 104100 195120 104120
rect 195380 104100 195620 104120
rect 195880 104100 196120 104120
rect 196380 104100 196620 104120
rect 196880 104100 197120 104120
rect 197380 104100 197620 104120
rect 197880 104100 198120 104120
rect 198380 104100 198620 104120
rect 198880 104100 199120 104120
rect 199380 104100 199620 104120
rect 199880 104100 200120 104120
rect 200380 104100 200620 104120
rect 200880 104100 201120 104120
rect 201380 104100 201620 104120
rect 201880 104100 202120 104120
rect 202380 104100 202620 104120
rect 202880 104100 203120 104120
rect 203380 104100 203620 104120
rect 203880 104100 204120 104120
rect 204380 104100 204620 104120
rect 204880 104100 205120 104120
rect 205380 104100 205620 104120
rect 205880 104100 206120 104120
rect 206380 104100 206620 104120
rect 206880 104100 207120 104120
rect 207380 104100 207620 104120
rect 207880 104100 208120 104120
rect 208380 104100 208620 104120
rect 208880 104100 209120 104120
rect 209380 104100 209620 104120
rect 209880 104100 210120 104120
rect 210380 104100 210620 104120
rect 210880 104100 211120 104120
rect 211380 104100 211620 104120
rect 211880 104100 212120 104120
rect 212380 104100 212620 104120
rect 212880 104100 213120 104120
rect 213380 104100 213620 104120
rect 213880 104100 214120 104120
rect 214380 104100 214620 104120
rect 214880 104100 215120 104120
rect 215380 104100 215620 104120
rect 215880 104100 216120 104120
rect 216380 104100 216620 104120
rect 216880 104100 217120 104120
rect 217380 104100 217620 104120
rect 217880 104100 218120 104120
rect 218380 104100 218620 104120
rect 218880 104100 219120 104120
rect 219380 104100 219620 104120
rect 219880 104100 220120 104120
rect 220380 104100 220620 104120
rect 220880 104100 221120 104120
rect 221380 104100 221620 104120
rect 221880 104100 222120 104120
rect 222380 104100 222620 104120
rect 222880 104100 223120 104120
rect 223380 104100 223620 104120
rect 223880 104100 224120 104120
rect 224380 104100 224620 104120
rect 224880 104100 225120 104120
rect 225380 104100 225620 104120
rect 225880 104100 226120 104120
rect 226380 104100 226620 104120
rect 226880 104100 227120 104120
rect 227380 104100 227620 104120
rect 227880 104100 228120 104120
rect 228380 104100 228620 104120
rect 228880 104100 229120 104120
rect 229380 104100 229620 104120
rect 229880 104100 230120 104120
rect 230380 104100 230620 104120
rect 230880 104100 231120 104120
rect 231380 104100 231620 104120
rect 231880 104100 232000 104120
rect 178000 104000 232000 104100
rect 178000 103900 188000 104000
rect 178000 103880 178120 103900
rect 178380 103880 178620 103900
rect 178880 103880 179120 103900
rect 179380 103880 179620 103900
rect 179880 103880 180120 103900
rect 180380 103880 180620 103900
rect 180880 103880 181120 103900
rect 181380 103880 181620 103900
rect 181880 103880 182120 103900
rect 182380 103880 182620 103900
rect 182880 103880 183120 103900
rect 183380 103880 183620 103900
rect 183880 103880 184120 103900
rect 184380 103880 184620 103900
rect 184880 103880 185120 103900
rect 185380 103880 185620 103900
rect 185880 103880 186120 103900
rect 186380 103880 186620 103900
rect 186880 103880 187120 103900
rect 187380 103880 187620 103900
rect 187880 103880 188000 103900
rect 178000 103620 178100 103880
rect 178400 103620 178600 103880
rect 178900 103620 179100 103880
rect 179400 103620 179600 103880
rect 179900 103620 180100 103880
rect 180400 103620 180600 103880
rect 180900 103620 181100 103880
rect 181400 103620 181600 103880
rect 181900 103620 182100 103880
rect 182400 103620 182600 103880
rect 182900 103620 183100 103880
rect 183400 103620 183600 103880
rect 183900 103620 184100 103880
rect 184400 103620 184600 103880
rect 184900 103620 185100 103880
rect 185400 103620 185600 103880
rect 185900 103620 186100 103880
rect 186400 103620 186600 103880
rect 186900 103620 187100 103880
rect 187400 103620 187600 103880
rect 187900 103620 188000 103880
rect 178000 103600 178120 103620
rect 178380 103600 178620 103620
rect 178880 103600 179120 103620
rect 179380 103600 179620 103620
rect 179880 103600 180120 103620
rect 180380 103600 180620 103620
rect 180880 103600 181120 103620
rect 181380 103600 181620 103620
rect 181880 103600 182120 103620
rect 182380 103600 182620 103620
rect 182880 103600 183120 103620
rect 183380 103600 183620 103620
rect 183880 103600 184120 103620
rect 184380 103600 184620 103620
rect 184880 103600 185120 103620
rect 185380 103600 185620 103620
rect 185880 103600 186120 103620
rect 186380 103600 186620 103620
rect 186880 103600 187120 103620
rect 187380 103600 187620 103620
rect 187880 103600 188000 103620
rect 178000 103400 188000 103600
rect 178000 103380 178120 103400
rect 178380 103380 178620 103400
rect 178880 103380 179120 103400
rect 179380 103380 179620 103400
rect 179880 103380 180120 103400
rect 180380 103380 180620 103400
rect 180880 103380 181120 103400
rect 181380 103380 181620 103400
rect 181880 103380 182120 103400
rect 182380 103380 182620 103400
rect 182880 103380 183120 103400
rect 183380 103380 183620 103400
rect 183880 103380 184120 103400
rect 184380 103380 184620 103400
rect 184880 103380 185120 103400
rect 185380 103380 185620 103400
rect 185880 103380 186120 103400
rect 186380 103380 186620 103400
rect 186880 103380 187120 103400
rect 187380 103380 187620 103400
rect 187880 103380 188000 103400
rect 178000 103120 178100 103380
rect 178400 103120 178600 103380
rect 178900 103120 179100 103380
rect 179400 103120 179600 103380
rect 179900 103120 180100 103380
rect 180400 103120 180600 103380
rect 180900 103120 181100 103380
rect 181400 103120 181600 103380
rect 181900 103120 182100 103380
rect 182400 103120 182600 103380
rect 182900 103120 183100 103380
rect 183400 103120 183600 103380
rect 183900 103120 184100 103380
rect 184400 103120 184600 103380
rect 184900 103120 185100 103380
rect 185400 103120 185600 103380
rect 185900 103120 186100 103380
rect 186400 103120 186600 103380
rect 186900 103120 187100 103380
rect 187400 103120 187600 103380
rect 187900 103120 188000 103380
rect 178000 103100 178120 103120
rect 178380 103100 178620 103120
rect 178880 103100 179120 103120
rect 179380 103100 179620 103120
rect 179880 103100 180120 103120
rect 180380 103100 180620 103120
rect 180880 103100 181120 103120
rect 181380 103100 181620 103120
rect 181880 103100 182120 103120
rect 182380 103100 182620 103120
rect 182880 103100 183120 103120
rect 183380 103100 183620 103120
rect 183880 103100 184120 103120
rect 184380 103100 184620 103120
rect 184880 103100 185120 103120
rect 185380 103100 185620 103120
rect 185880 103100 186120 103120
rect 186380 103100 186620 103120
rect 186880 103100 187120 103120
rect 187380 103100 187620 103120
rect 187880 103100 188000 103120
rect 178000 102900 188000 103100
rect 178000 102880 178120 102900
rect 178380 102880 178620 102900
rect 178880 102880 179120 102900
rect 179380 102880 179620 102900
rect 179880 102880 180120 102900
rect 180380 102880 180620 102900
rect 180880 102880 181120 102900
rect 181380 102880 181620 102900
rect 181880 102880 182120 102900
rect 182380 102880 182620 102900
rect 182880 102880 183120 102900
rect 183380 102880 183620 102900
rect 183880 102880 184120 102900
rect 184380 102880 184620 102900
rect 184880 102880 185120 102900
rect 185380 102880 185620 102900
rect 185880 102880 186120 102900
rect 186380 102880 186620 102900
rect 186880 102880 187120 102900
rect 187380 102880 187620 102900
rect 187880 102880 188000 102900
rect 178000 102620 178100 102880
rect 178400 102620 178600 102880
rect 178900 102620 179100 102880
rect 179400 102620 179600 102880
rect 179900 102620 180100 102880
rect 180400 102620 180600 102880
rect 180900 102620 181100 102880
rect 181400 102620 181600 102880
rect 181900 102620 182100 102880
rect 182400 102620 182600 102880
rect 182900 102620 183100 102880
rect 183400 102620 183600 102880
rect 183900 102620 184100 102880
rect 184400 102620 184600 102880
rect 184900 102620 185100 102880
rect 185400 102620 185600 102880
rect 185900 102620 186100 102880
rect 186400 102620 186600 102880
rect 186900 102620 187100 102880
rect 187400 102620 187600 102880
rect 187900 102620 188000 102880
rect 178000 102600 178120 102620
rect 178380 102600 178620 102620
rect 178880 102600 179120 102620
rect 179380 102600 179620 102620
rect 179880 102600 180120 102620
rect 180380 102600 180620 102620
rect 180880 102600 181120 102620
rect 181380 102600 181620 102620
rect 181880 102600 182120 102620
rect 182380 102600 182620 102620
rect 182880 102600 183120 102620
rect 183380 102600 183620 102620
rect 183880 102600 184120 102620
rect 184380 102600 184620 102620
rect 184880 102600 185120 102620
rect 185380 102600 185620 102620
rect 185880 102600 186120 102620
rect 186380 102600 186620 102620
rect 186880 102600 187120 102620
rect 187380 102600 187620 102620
rect 187880 102600 188000 102620
rect 178000 102400 188000 102600
rect 178000 102380 178120 102400
rect 178380 102380 178620 102400
rect 178880 102380 179120 102400
rect 179380 102380 179620 102400
rect 179880 102380 180120 102400
rect 180380 102380 180620 102400
rect 180880 102380 181120 102400
rect 181380 102380 181620 102400
rect 181880 102380 182120 102400
rect 182380 102380 182620 102400
rect 182880 102380 183120 102400
rect 183380 102380 183620 102400
rect 183880 102380 184120 102400
rect 184380 102380 184620 102400
rect 184880 102380 185120 102400
rect 185380 102380 185620 102400
rect 185880 102380 186120 102400
rect 186380 102380 186620 102400
rect 186880 102380 187120 102400
rect 187380 102380 187620 102400
rect 187880 102380 188000 102400
rect 178000 102120 178100 102380
rect 178400 102120 178600 102380
rect 178900 102120 179100 102380
rect 179400 102120 179600 102380
rect 179900 102120 180100 102380
rect 180400 102120 180600 102380
rect 180900 102120 181100 102380
rect 181400 102120 181600 102380
rect 181900 102120 182100 102380
rect 182400 102120 182600 102380
rect 182900 102120 183100 102380
rect 183400 102120 183600 102380
rect 183900 102120 184100 102380
rect 184400 102120 184600 102380
rect 184900 102120 185100 102380
rect 185400 102120 185600 102380
rect 185900 102120 186100 102380
rect 186400 102120 186600 102380
rect 186900 102120 187100 102380
rect 187400 102120 187600 102380
rect 187900 102120 188000 102380
rect 178000 102100 178120 102120
rect 178380 102100 178620 102120
rect 178880 102100 179120 102120
rect 179380 102100 179620 102120
rect 179880 102100 180120 102120
rect 180380 102100 180620 102120
rect 180880 102100 181120 102120
rect 181380 102100 181620 102120
rect 181880 102100 182120 102120
rect 182380 102100 182620 102120
rect 182880 102100 183120 102120
rect 183380 102100 183620 102120
rect 183880 102100 184120 102120
rect 184380 102100 184620 102120
rect 184880 102100 185120 102120
rect 185380 102100 185620 102120
rect 185880 102100 186120 102120
rect 186380 102100 186620 102120
rect 186880 102100 187120 102120
rect 187380 102100 187620 102120
rect 187880 102100 188000 102120
rect 178000 102000 188000 102100
rect 196000 103980 208000 104000
rect 196000 103910 196150 103980
rect 196350 103910 196650 103980
rect 196850 103910 197150 103980
rect 197350 103910 197650 103980
rect 197850 103910 198150 103980
rect 198350 103910 198650 103980
rect 198850 103910 199150 103980
rect 199350 103910 199650 103980
rect 199850 103910 200150 103980
rect 200350 103910 200650 103980
rect 200850 103910 201150 103980
rect 201350 103910 201650 103980
rect 201850 103910 202150 103980
rect 202350 103910 202650 103980
rect 202850 103910 203150 103980
rect 203350 103910 203650 103980
rect 203850 103910 204150 103980
rect 204350 103910 204650 103980
rect 204850 103910 205150 103980
rect 205350 103910 205650 103980
rect 205850 103910 206150 103980
rect 206350 103910 206650 103980
rect 206850 103910 207150 103980
rect 207350 103910 207650 103980
rect 207850 103910 208000 103980
rect 196000 103900 208000 103910
rect 196000 103880 196120 103900
rect 196380 103880 196620 103900
rect 196880 103880 197120 103900
rect 197380 103880 197620 103900
rect 197880 103880 198120 103900
rect 198380 103880 198620 103900
rect 198880 103880 199120 103900
rect 199380 103880 199620 103900
rect 199880 103880 200120 103900
rect 200380 103880 200620 103900
rect 200880 103880 201120 103900
rect 201380 103880 201620 103900
rect 201880 103880 202120 103900
rect 202380 103880 202620 103900
rect 202880 103880 203120 103900
rect 203380 103880 203620 103900
rect 203880 103880 204120 103900
rect 204380 103880 204620 103900
rect 204880 103880 205120 103900
rect 205380 103880 205620 103900
rect 205880 103880 206120 103900
rect 206380 103880 206620 103900
rect 206880 103880 207120 103900
rect 207380 103880 207620 103900
rect 207880 103880 208000 103900
rect 196000 103850 196100 103880
rect 196000 103650 196020 103850
rect 196090 103650 196100 103850
rect 196000 103620 196100 103650
rect 196400 103850 196600 103880
rect 196400 103650 196410 103850
rect 196480 103650 196520 103850
rect 196590 103650 196600 103850
rect 196400 103620 196600 103650
rect 196900 103850 197100 103880
rect 196900 103650 196910 103850
rect 196980 103650 197020 103850
rect 197090 103650 197100 103850
rect 196900 103620 197100 103650
rect 197400 103850 197600 103880
rect 197400 103650 197410 103850
rect 197480 103650 197520 103850
rect 197590 103650 197600 103850
rect 197400 103620 197600 103650
rect 197900 103850 198100 103880
rect 197900 103650 197910 103850
rect 197980 103650 198020 103850
rect 198090 103650 198100 103850
rect 197900 103620 198100 103650
rect 198400 103850 198600 103880
rect 198400 103650 198410 103850
rect 198480 103650 198520 103850
rect 198590 103650 198600 103850
rect 198400 103620 198600 103650
rect 198900 103850 199100 103880
rect 198900 103650 198910 103850
rect 198980 103650 199020 103850
rect 199090 103650 199100 103850
rect 198900 103620 199100 103650
rect 199400 103850 199600 103880
rect 199400 103650 199410 103850
rect 199480 103650 199520 103850
rect 199590 103650 199600 103850
rect 199400 103620 199600 103650
rect 199900 103850 200100 103880
rect 199900 103650 199910 103850
rect 199980 103650 200020 103850
rect 200090 103650 200100 103850
rect 199900 103620 200100 103650
rect 200400 103850 200600 103880
rect 200400 103650 200410 103850
rect 200480 103650 200520 103850
rect 200590 103650 200600 103850
rect 200400 103620 200600 103650
rect 200900 103850 201100 103880
rect 200900 103650 200910 103850
rect 200980 103650 201020 103850
rect 201090 103650 201100 103850
rect 200900 103620 201100 103650
rect 201400 103850 201600 103880
rect 201400 103650 201410 103850
rect 201480 103650 201520 103850
rect 201590 103650 201600 103850
rect 201400 103620 201600 103650
rect 201900 103850 202100 103880
rect 201900 103650 201910 103850
rect 201980 103650 202020 103850
rect 202090 103650 202100 103850
rect 201900 103620 202100 103650
rect 202400 103850 202600 103880
rect 202400 103650 202410 103850
rect 202480 103650 202520 103850
rect 202590 103650 202600 103850
rect 202400 103620 202600 103650
rect 202900 103850 203100 103880
rect 202900 103650 202910 103850
rect 202980 103650 203020 103850
rect 203090 103650 203100 103850
rect 202900 103620 203100 103650
rect 203400 103850 203600 103880
rect 203400 103650 203410 103850
rect 203480 103650 203520 103850
rect 203590 103650 203600 103850
rect 203400 103620 203600 103650
rect 203900 103850 204100 103880
rect 203900 103650 203910 103850
rect 203980 103650 204020 103850
rect 204090 103650 204100 103850
rect 203900 103620 204100 103650
rect 204400 103850 204600 103880
rect 204400 103650 204410 103850
rect 204480 103650 204520 103850
rect 204590 103650 204600 103850
rect 204400 103620 204600 103650
rect 204900 103850 205100 103880
rect 204900 103650 204910 103850
rect 204980 103650 205020 103850
rect 205090 103650 205100 103850
rect 204900 103620 205100 103650
rect 205400 103850 205600 103880
rect 205400 103650 205410 103850
rect 205480 103650 205520 103850
rect 205590 103650 205600 103850
rect 205400 103620 205600 103650
rect 205900 103850 206100 103880
rect 205900 103650 205910 103850
rect 205980 103650 206020 103850
rect 206090 103650 206100 103850
rect 205900 103620 206100 103650
rect 206400 103850 206600 103880
rect 206400 103650 206410 103850
rect 206480 103650 206520 103850
rect 206590 103650 206600 103850
rect 206400 103620 206600 103650
rect 206900 103850 207100 103880
rect 206900 103650 206910 103850
rect 206980 103650 207020 103850
rect 207090 103650 207100 103850
rect 206900 103620 207100 103650
rect 207400 103850 207600 103880
rect 207400 103650 207410 103850
rect 207480 103650 207520 103850
rect 207590 103650 207600 103850
rect 207400 103620 207600 103650
rect 207900 103850 208000 103880
rect 207900 103650 207910 103850
rect 207980 103650 208000 103850
rect 207900 103620 208000 103650
rect 196000 103600 196120 103620
rect 196380 103600 196620 103620
rect 196880 103600 197120 103620
rect 197380 103600 197620 103620
rect 197880 103600 198120 103620
rect 198380 103600 198620 103620
rect 198880 103600 199120 103620
rect 199380 103600 199620 103620
rect 199880 103600 200120 103620
rect 200380 103600 200620 103620
rect 200880 103600 201120 103620
rect 201380 103600 201620 103620
rect 201880 103600 202120 103620
rect 202380 103600 202620 103620
rect 202880 103600 203120 103620
rect 203380 103600 203620 103620
rect 203880 103600 204120 103620
rect 204380 103600 204620 103620
rect 204880 103600 205120 103620
rect 205380 103600 205620 103620
rect 205880 103600 206120 103620
rect 206380 103600 206620 103620
rect 206880 103600 207120 103620
rect 207380 103600 207620 103620
rect 207880 103600 208000 103620
rect 196000 103590 208000 103600
rect 196000 103520 196150 103590
rect 196350 103520 196650 103590
rect 196850 103520 197150 103590
rect 197350 103520 197650 103590
rect 197850 103520 198150 103590
rect 198350 103520 198650 103590
rect 198850 103520 199150 103590
rect 199350 103520 199650 103590
rect 199850 103520 200150 103590
rect 200350 103520 200650 103590
rect 200850 103520 201150 103590
rect 201350 103520 201650 103590
rect 201850 103520 202150 103590
rect 202350 103520 202650 103590
rect 202850 103520 203150 103590
rect 203350 103520 203650 103590
rect 203850 103520 204150 103590
rect 204350 103520 204650 103590
rect 204850 103520 205150 103590
rect 205350 103520 205650 103590
rect 205850 103520 206150 103590
rect 206350 103520 206650 103590
rect 206850 103520 207150 103590
rect 207350 103520 207650 103590
rect 207850 103520 208000 103590
rect 196000 103480 208000 103520
rect 196000 103410 196150 103480
rect 196350 103410 196650 103480
rect 196850 103410 197150 103480
rect 197350 103410 197650 103480
rect 197850 103410 198150 103480
rect 198350 103410 198650 103480
rect 198850 103410 199150 103480
rect 199350 103410 199650 103480
rect 199850 103410 200150 103480
rect 200350 103410 200650 103480
rect 200850 103410 201150 103480
rect 201350 103410 201650 103480
rect 201850 103410 202150 103480
rect 202350 103410 202650 103480
rect 202850 103410 203150 103480
rect 203350 103410 203650 103480
rect 203850 103410 204150 103480
rect 204350 103410 204650 103480
rect 204850 103410 205150 103480
rect 205350 103410 205650 103480
rect 205850 103410 206150 103480
rect 206350 103410 206650 103480
rect 206850 103410 207150 103480
rect 207350 103410 207650 103480
rect 207850 103410 208000 103480
rect 196000 103400 208000 103410
rect 196000 103380 196120 103400
rect 196380 103380 196620 103400
rect 196880 103380 197120 103400
rect 197380 103380 197620 103400
rect 197880 103380 198120 103400
rect 198380 103380 198620 103400
rect 198880 103380 199120 103400
rect 199380 103380 199620 103400
rect 199880 103380 200120 103400
rect 200380 103380 200620 103400
rect 200880 103380 201120 103400
rect 201380 103380 201620 103400
rect 201880 103380 202120 103400
rect 202380 103380 202620 103400
rect 202880 103380 203120 103400
rect 203380 103380 203620 103400
rect 203880 103380 204120 103400
rect 204380 103380 204620 103400
rect 204880 103380 205120 103400
rect 205380 103380 205620 103400
rect 205880 103380 206120 103400
rect 206380 103380 206620 103400
rect 206880 103380 207120 103400
rect 207380 103380 207620 103400
rect 207880 103380 208000 103400
rect 196000 103350 196100 103380
rect 196000 103150 196020 103350
rect 196090 103150 196100 103350
rect 196000 103120 196100 103150
rect 196400 103350 196600 103380
rect 196400 103150 196410 103350
rect 196480 103150 196520 103350
rect 196590 103150 196600 103350
rect 196400 103120 196600 103150
rect 196900 103350 197100 103380
rect 196900 103150 196910 103350
rect 196980 103150 197020 103350
rect 197090 103150 197100 103350
rect 196900 103120 197100 103150
rect 197400 103350 197600 103380
rect 197400 103150 197410 103350
rect 197480 103150 197520 103350
rect 197590 103150 197600 103350
rect 197400 103120 197600 103150
rect 197900 103350 198100 103380
rect 197900 103150 197910 103350
rect 197980 103150 198020 103350
rect 198090 103150 198100 103350
rect 197900 103120 198100 103150
rect 198400 103350 198600 103380
rect 198400 103150 198410 103350
rect 198480 103150 198520 103350
rect 198590 103150 198600 103350
rect 198400 103120 198600 103150
rect 198900 103350 199100 103380
rect 198900 103150 198910 103350
rect 198980 103150 199020 103350
rect 199090 103150 199100 103350
rect 198900 103120 199100 103150
rect 199400 103350 199600 103380
rect 199400 103150 199410 103350
rect 199480 103150 199520 103350
rect 199590 103150 199600 103350
rect 199400 103120 199600 103150
rect 199900 103350 200100 103380
rect 199900 103150 199910 103350
rect 199980 103150 200020 103350
rect 200090 103150 200100 103350
rect 199900 103120 200100 103150
rect 200400 103350 200600 103380
rect 200400 103150 200410 103350
rect 200480 103150 200520 103350
rect 200590 103150 200600 103350
rect 200400 103120 200600 103150
rect 200900 103350 201100 103380
rect 200900 103150 200910 103350
rect 200980 103150 201020 103350
rect 201090 103150 201100 103350
rect 200900 103120 201100 103150
rect 201400 103350 201600 103380
rect 201400 103150 201410 103350
rect 201480 103150 201520 103350
rect 201590 103150 201600 103350
rect 201400 103120 201600 103150
rect 201900 103350 202100 103380
rect 201900 103150 201910 103350
rect 201980 103150 202020 103350
rect 202090 103150 202100 103350
rect 201900 103120 202100 103150
rect 202400 103350 202600 103380
rect 202400 103150 202410 103350
rect 202480 103150 202520 103350
rect 202590 103150 202600 103350
rect 202400 103120 202600 103150
rect 202900 103350 203100 103380
rect 202900 103150 202910 103350
rect 202980 103150 203020 103350
rect 203090 103150 203100 103350
rect 202900 103120 203100 103150
rect 203400 103350 203600 103380
rect 203400 103150 203410 103350
rect 203480 103150 203520 103350
rect 203590 103150 203600 103350
rect 203400 103120 203600 103150
rect 203900 103350 204100 103380
rect 203900 103150 203910 103350
rect 203980 103150 204020 103350
rect 204090 103150 204100 103350
rect 203900 103120 204100 103150
rect 204400 103350 204600 103380
rect 204400 103150 204410 103350
rect 204480 103150 204520 103350
rect 204590 103150 204600 103350
rect 204400 103120 204600 103150
rect 204900 103350 205100 103380
rect 204900 103150 204910 103350
rect 204980 103150 205020 103350
rect 205090 103150 205100 103350
rect 204900 103120 205100 103150
rect 205400 103350 205600 103380
rect 205400 103150 205410 103350
rect 205480 103150 205520 103350
rect 205590 103150 205600 103350
rect 205400 103120 205600 103150
rect 205900 103350 206100 103380
rect 205900 103150 205910 103350
rect 205980 103150 206020 103350
rect 206090 103150 206100 103350
rect 205900 103120 206100 103150
rect 206400 103350 206600 103380
rect 206400 103150 206410 103350
rect 206480 103150 206520 103350
rect 206590 103150 206600 103350
rect 206400 103120 206600 103150
rect 206900 103350 207100 103380
rect 206900 103150 206910 103350
rect 206980 103150 207020 103350
rect 207090 103150 207100 103350
rect 206900 103120 207100 103150
rect 207400 103350 207600 103380
rect 207400 103150 207410 103350
rect 207480 103150 207520 103350
rect 207590 103150 207600 103350
rect 207400 103120 207600 103150
rect 207900 103350 208000 103380
rect 207900 103150 207910 103350
rect 207980 103150 208000 103350
rect 207900 103120 208000 103150
rect 196000 103100 196120 103120
rect 196380 103100 196620 103120
rect 196880 103100 197120 103120
rect 197380 103100 197620 103120
rect 197880 103100 198120 103120
rect 198380 103100 198620 103120
rect 198880 103100 199120 103120
rect 199380 103100 199620 103120
rect 199880 103100 200120 103120
rect 200380 103100 200620 103120
rect 200880 103100 201120 103120
rect 201380 103100 201620 103120
rect 201880 103100 202120 103120
rect 202380 103100 202620 103120
rect 202880 103100 203120 103120
rect 203380 103100 203620 103120
rect 203880 103100 204120 103120
rect 204380 103100 204620 103120
rect 204880 103100 205120 103120
rect 205380 103100 205620 103120
rect 205880 103100 206120 103120
rect 206380 103100 206620 103120
rect 206880 103100 207120 103120
rect 207380 103100 207620 103120
rect 207880 103100 208000 103120
rect 196000 103090 208000 103100
rect 196000 103020 196150 103090
rect 196350 103020 196650 103090
rect 196850 103020 197150 103090
rect 197350 103020 197650 103090
rect 197850 103020 198150 103090
rect 198350 103020 198650 103090
rect 198850 103020 199150 103090
rect 199350 103020 199650 103090
rect 199850 103020 200150 103090
rect 200350 103020 200650 103090
rect 200850 103020 201150 103090
rect 201350 103020 201650 103090
rect 201850 103020 202150 103090
rect 202350 103020 202650 103090
rect 202850 103020 203150 103090
rect 203350 103020 203650 103090
rect 203850 103020 204150 103090
rect 204350 103020 204650 103090
rect 204850 103020 205150 103090
rect 205350 103020 205650 103090
rect 205850 103020 206150 103090
rect 206350 103020 206650 103090
rect 206850 103020 207150 103090
rect 207350 103020 207650 103090
rect 207850 103020 208000 103090
rect 196000 102980 208000 103020
rect 196000 102910 196150 102980
rect 196350 102910 196650 102980
rect 196850 102910 197150 102980
rect 197350 102910 197650 102980
rect 197850 102910 198150 102980
rect 198350 102910 198650 102980
rect 198850 102910 199150 102980
rect 199350 102910 199650 102980
rect 199850 102910 200150 102980
rect 200350 102910 200650 102980
rect 200850 102910 201150 102980
rect 201350 102910 201650 102980
rect 201850 102910 202150 102980
rect 202350 102910 202650 102980
rect 202850 102910 203150 102980
rect 203350 102910 203650 102980
rect 203850 102910 204150 102980
rect 204350 102910 204650 102980
rect 204850 102910 205150 102980
rect 205350 102910 205650 102980
rect 205850 102910 206150 102980
rect 206350 102910 206650 102980
rect 206850 102910 207150 102980
rect 207350 102910 207650 102980
rect 207850 102910 208000 102980
rect 196000 102900 208000 102910
rect 196000 102880 196120 102900
rect 196380 102880 196620 102900
rect 196880 102880 197120 102900
rect 197380 102880 197620 102900
rect 197880 102880 198120 102900
rect 198380 102880 198620 102900
rect 198880 102880 199120 102900
rect 199380 102880 199620 102900
rect 199880 102880 200120 102900
rect 200380 102880 200620 102900
rect 200880 102880 201120 102900
rect 201380 102880 201620 102900
rect 201880 102880 202120 102900
rect 202380 102880 202620 102900
rect 202880 102880 203120 102900
rect 203380 102880 203620 102900
rect 203880 102880 204120 102900
rect 204380 102880 204620 102900
rect 204880 102880 205120 102900
rect 205380 102880 205620 102900
rect 205880 102880 206120 102900
rect 206380 102880 206620 102900
rect 206880 102880 207120 102900
rect 207380 102880 207620 102900
rect 207880 102880 208000 102900
rect 196000 102850 196100 102880
rect 196000 102650 196020 102850
rect 196090 102650 196100 102850
rect 196000 102620 196100 102650
rect 196400 102850 196600 102880
rect 196400 102650 196410 102850
rect 196480 102650 196520 102850
rect 196590 102650 196600 102850
rect 196400 102620 196600 102650
rect 196900 102850 197100 102880
rect 196900 102650 196910 102850
rect 196980 102650 197020 102850
rect 197090 102650 197100 102850
rect 196900 102620 197100 102650
rect 197400 102850 197600 102880
rect 197400 102650 197410 102850
rect 197480 102650 197520 102850
rect 197590 102650 197600 102850
rect 197400 102620 197600 102650
rect 197900 102850 198100 102880
rect 197900 102650 197910 102850
rect 197980 102650 198020 102850
rect 198090 102650 198100 102850
rect 197900 102620 198100 102650
rect 198400 102850 198600 102880
rect 198400 102650 198410 102850
rect 198480 102650 198520 102850
rect 198590 102650 198600 102850
rect 198400 102620 198600 102650
rect 198900 102850 199100 102880
rect 198900 102650 198910 102850
rect 198980 102650 199020 102850
rect 199090 102650 199100 102850
rect 198900 102620 199100 102650
rect 199400 102850 199600 102880
rect 199400 102650 199410 102850
rect 199480 102650 199520 102850
rect 199590 102650 199600 102850
rect 199400 102620 199600 102650
rect 199900 102850 200100 102880
rect 199900 102650 199910 102850
rect 199980 102650 200020 102850
rect 200090 102650 200100 102850
rect 199900 102620 200100 102650
rect 200400 102850 200600 102880
rect 200400 102650 200410 102850
rect 200480 102650 200520 102850
rect 200590 102650 200600 102850
rect 200400 102620 200600 102650
rect 200900 102850 201100 102880
rect 200900 102650 200910 102850
rect 200980 102650 201020 102850
rect 201090 102650 201100 102850
rect 200900 102620 201100 102650
rect 201400 102850 201600 102880
rect 201400 102650 201410 102850
rect 201480 102650 201520 102850
rect 201590 102650 201600 102850
rect 201400 102620 201600 102650
rect 201900 102850 202100 102880
rect 201900 102650 201910 102850
rect 201980 102650 202020 102850
rect 202090 102650 202100 102850
rect 201900 102620 202100 102650
rect 202400 102850 202600 102880
rect 202400 102650 202410 102850
rect 202480 102650 202520 102850
rect 202590 102650 202600 102850
rect 202400 102620 202600 102650
rect 202900 102850 203100 102880
rect 202900 102650 202910 102850
rect 202980 102650 203020 102850
rect 203090 102650 203100 102850
rect 202900 102620 203100 102650
rect 203400 102850 203600 102880
rect 203400 102650 203410 102850
rect 203480 102650 203520 102850
rect 203590 102650 203600 102850
rect 203400 102620 203600 102650
rect 203900 102850 204100 102880
rect 203900 102650 203910 102850
rect 203980 102650 204020 102850
rect 204090 102650 204100 102850
rect 203900 102620 204100 102650
rect 204400 102850 204600 102880
rect 204400 102650 204410 102850
rect 204480 102650 204520 102850
rect 204590 102650 204600 102850
rect 204400 102620 204600 102650
rect 204900 102850 205100 102880
rect 204900 102650 204910 102850
rect 204980 102650 205020 102850
rect 205090 102650 205100 102850
rect 204900 102620 205100 102650
rect 205400 102850 205600 102880
rect 205400 102650 205410 102850
rect 205480 102650 205520 102850
rect 205590 102650 205600 102850
rect 205400 102620 205600 102650
rect 205900 102850 206100 102880
rect 205900 102650 205910 102850
rect 205980 102650 206020 102850
rect 206090 102650 206100 102850
rect 205900 102620 206100 102650
rect 206400 102850 206600 102880
rect 206400 102650 206410 102850
rect 206480 102650 206520 102850
rect 206590 102650 206600 102850
rect 206400 102620 206600 102650
rect 206900 102850 207100 102880
rect 206900 102650 206910 102850
rect 206980 102650 207020 102850
rect 207090 102650 207100 102850
rect 206900 102620 207100 102650
rect 207400 102850 207600 102880
rect 207400 102650 207410 102850
rect 207480 102650 207520 102850
rect 207590 102650 207600 102850
rect 207400 102620 207600 102650
rect 207900 102850 208000 102880
rect 207900 102650 207910 102850
rect 207980 102650 208000 102850
rect 207900 102620 208000 102650
rect 196000 102600 196120 102620
rect 196380 102600 196620 102620
rect 196880 102600 197120 102620
rect 197380 102600 197620 102620
rect 197880 102600 198120 102620
rect 198380 102600 198620 102620
rect 198880 102600 199120 102620
rect 199380 102600 199620 102620
rect 199880 102600 200120 102620
rect 200380 102600 200620 102620
rect 200880 102600 201120 102620
rect 201380 102600 201620 102620
rect 201880 102600 202120 102620
rect 202380 102600 202620 102620
rect 202880 102600 203120 102620
rect 203380 102600 203620 102620
rect 203880 102600 204120 102620
rect 204380 102600 204620 102620
rect 204880 102600 205120 102620
rect 205380 102600 205620 102620
rect 205880 102600 206120 102620
rect 206380 102600 206620 102620
rect 206880 102600 207120 102620
rect 207380 102600 207620 102620
rect 207880 102600 208000 102620
rect 196000 102590 208000 102600
rect 196000 102520 196150 102590
rect 196350 102520 196650 102590
rect 196850 102520 197150 102590
rect 197350 102520 197650 102590
rect 197850 102520 198150 102590
rect 198350 102520 198650 102590
rect 198850 102520 199150 102590
rect 199350 102520 199650 102590
rect 199850 102520 200150 102590
rect 200350 102520 200650 102590
rect 200850 102520 201150 102590
rect 201350 102520 201650 102590
rect 201850 102520 202150 102590
rect 202350 102520 202650 102590
rect 202850 102520 203150 102590
rect 203350 102520 203650 102590
rect 203850 102520 204150 102590
rect 204350 102520 204650 102590
rect 204850 102520 205150 102590
rect 205350 102520 205650 102590
rect 205850 102520 206150 102590
rect 206350 102520 206650 102590
rect 206850 102520 207150 102590
rect 207350 102520 207650 102590
rect 207850 102520 208000 102590
rect 196000 102480 208000 102520
rect 196000 102410 196150 102480
rect 196350 102410 196650 102480
rect 196850 102410 197150 102480
rect 197350 102410 197650 102480
rect 197850 102410 198150 102480
rect 198350 102410 198650 102480
rect 198850 102410 199150 102480
rect 199350 102410 199650 102480
rect 199850 102410 200150 102480
rect 200350 102410 200650 102480
rect 200850 102410 201150 102480
rect 201350 102410 201650 102480
rect 201850 102410 202150 102480
rect 202350 102410 202650 102480
rect 202850 102410 203150 102480
rect 203350 102410 203650 102480
rect 203850 102410 204150 102480
rect 204350 102410 204650 102480
rect 204850 102410 205150 102480
rect 205350 102410 205650 102480
rect 205850 102410 206150 102480
rect 206350 102410 206650 102480
rect 206850 102410 207150 102480
rect 207350 102410 207650 102480
rect 207850 102410 208000 102480
rect 196000 102400 208000 102410
rect 196000 102380 196120 102400
rect 196380 102380 196620 102400
rect 196880 102380 197120 102400
rect 197380 102380 197620 102400
rect 197880 102380 198120 102400
rect 198380 102380 198620 102400
rect 198880 102380 199120 102400
rect 199380 102380 199620 102400
rect 199880 102380 200120 102400
rect 200380 102380 200620 102400
rect 200880 102380 201120 102400
rect 201380 102380 201620 102400
rect 201880 102380 202120 102400
rect 202380 102380 202620 102400
rect 202880 102380 203120 102400
rect 203380 102380 203620 102400
rect 203880 102380 204120 102400
rect 204380 102380 204620 102400
rect 204880 102380 205120 102400
rect 205380 102380 205620 102400
rect 205880 102380 206120 102400
rect 206380 102380 206620 102400
rect 206880 102380 207120 102400
rect 207380 102380 207620 102400
rect 207880 102380 208000 102400
rect 196000 102350 196100 102380
rect 196000 102150 196020 102350
rect 196090 102150 196100 102350
rect 196000 102120 196100 102150
rect 196400 102350 196600 102380
rect 196400 102150 196410 102350
rect 196480 102150 196520 102350
rect 196590 102150 196600 102350
rect 196400 102120 196600 102150
rect 196900 102350 197100 102380
rect 196900 102150 196910 102350
rect 196980 102150 197020 102350
rect 197090 102150 197100 102350
rect 196900 102120 197100 102150
rect 197400 102350 197600 102380
rect 197400 102150 197410 102350
rect 197480 102150 197520 102350
rect 197590 102150 197600 102350
rect 197400 102120 197600 102150
rect 197900 102350 198100 102380
rect 197900 102150 197910 102350
rect 197980 102150 198020 102350
rect 198090 102150 198100 102350
rect 197900 102120 198100 102150
rect 198400 102350 198600 102380
rect 198400 102150 198410 102350
rect 198480 102150 198520 102350
rect 198590 102150 198600 102350
rect 198400 102120 198600 102150
rect 198900 102350 199100 102380
rect 198900 102150 198910 102350
rect 198980 102150 199020 102350
rect 199090 102150 199100 102350
rect 198900 102120 199100 102150
rect 199400 102350 199600 102380
rect 199400 102150 199410 102350
rect 199480 102150 199520 102350
rect 199590 102150 199600 102350
rect 199400 102120 199600 102150
rect 199900 102350 200100 102380
rect 199900 102150 199910 102350
rect 199980 102150 200020 102350
rect 200090 102150 200100 102350
rect 199900 102120 200100 102150
rect 200400 102350 200600 102380
rect 200400 102150 200410 102350
rect 200480 102150 200520 102350
rect 200590 102150 200600 102350
rect 200400 102120 200600 102150
rect 200900 102350 201100 102380
rect 200900 102150 200910 102350
rect 200980 102150 201020 102350
rect 201090 102150 201100 102350
rect 200900 102120 201100 102150
rect 201400 102350 201600 102380
rect 201400 102150 201410 102350
rect 201480 102150 201520 102350
rect 201590 102150 201600 102350
rect 201400 102120 201600 102150
rect 201900 102350 202100 102380
rect 201900 102150 201910 102350
rect 201980 102150 202020 102350
rect 202090 102150 202100 102350
rect 201900 102120 202100 102150
rect 202400 102350 202600 102380
rect 202400 102150 202410 102350
rect 202480 102150 202520 102350
rect 202590 102150 202600 102350
rect 202400 102120 202600 102150
rect 202900 102350 203100 102380
rect 202900 102150 202910 102350
rect 202980 102150 203020 102350
rect 203090 102150 203100 102350
rect 202900 102120 203100 102150
rect 203400 102350 203600 102380
rect 203400 102150 203410 102350
rect 203480 102150 203520 102350
rect 203590 102150 203600 102350
rect 203400 102120 203600 102150
rect 203900 102350 204100 102380
rect 203900 102150 203910 102350
rect 203980 102150 204020 102350
rect 204090 102150 204100 102350
rect 203900 102120 204100 102150
rect 204400 102350 204600 102380
rect 204400 102150 204410 102350
rect 204480 102150 204520 102350
rect 204590 102150 204600 102350
rect 204400 102120 204600 102150
rect 204900 102350 205100 102380
rect 204900 102150 204910 102350
rect 204980 102150 205020 102350
rect 205090 102150 205100 102350
rect 204900 102120 205100 102150
rect 205400 102350 205600 102380
rect 205400 102150 205410 102350
rect 205480 102150 205520 102350
rect 205590 102150 205600 102350
rect 205400 102120 205600 102150
rect 205900 102350 206100 102380
rect 205900 102150 205910 102350
rect 205980 102150 206020 102350
rect 206090 102150 206100 102350
rect 205900 102120 206100 102150
rect 206400 102350 206600 102380
rect 206400 102150 206410 102350
rect 206480 102150 206520 102350
rect 206590 102150 206600 102350
rect 206400 102120 206600 102150
rect 206900 102350 207100 102380
rect 206900 102150 206910 102350
rect 206980 102150 207020 102350
rect 207090 102150 207100 102350
rect 206900 102120 207100 102150
rect 207400 102350 207600 102380
rect 207400 102150 207410 102350
rect 207480 102150 207520 102350
rect 207590 102150 207600 102350
rect 207400 102120 207600 102150
rect 207900 102350 208000 102380
rect 207900 102150 207910 102350
rect 207980 102150 208000 102350
rect 207900 102120 208000 102150
rect 196000 102100 196120 102120
rect 196380 102100 196620 102120
rect 196880 102100 197120 102120
rect 197380 102100 197620 102120
rect 197880 102100 198120 102120
rect 198380 102100 198620 102120
rect 198880 102100 199120 102120
rect 199380 102100 199620 102120
rect 199880 102100 200120 102120
rect 200380 102100 200620 102120
rect 200880 102100 201120 102120
rect 201380 102100 201620 102120
rect 201880 102100 202120 102120
rect 202380 102100 202620 102120
rect 202880 102100 203120 102120
rect 203380 102100 203620 102120
rect 203880 102100 204120 102120
rect 204380 102100 204620 102120
rect 204880 102100 205120 102120
rect 205380 102100 205620 102120
rect 205880 102100 206120 102120
rect 206380 102100 206620 102120
rect 206880 102100 207120 102120
rect 207380 102100 207620 102120
rect 207880 102100 208000 102120
rect 196000 102090 208000 102100
rect 196000 102020 196150 102090
rect 196350 102020 196650 102090
rect 196850 102020 197150 102090
rect 197350 102020 197650 102090
rect 197850 102020 198150 102090
rect 198350 102020 198650 102090
rect 198850 102020 199150 102090
rect 199350 102020 199650 102090
rect 199850 102020 200150 102090
rect 200350 102020 200650 102090
rect 200850 102020 201150 102090
rect 201350 102020 201650 102090
rect 201850 102020 202150 102090
rect 202350 102020 202650 102090
rect 202850 102020 203150 102090
rect 203350 102020 203650 102090
rect 203850 102020 204150 102090
rect 204350 102020 204650 102090
rect 204850 102020 205150 102090
rect 205350 102020 205650 102090
rect 205850 102020 206150 102090
rect 206350 102020 206650 102090
rect 206850 102020 207150 102090
rect 207350 102020 207650 102090
rect 207850 102020 208000 102090
rect 196000 101980 208000 102020
rect 196000 101910 196150 101980
rect 196350 101910 196650 101980
rect 196850 101910 197150 101980
rect 197350 101910 197650 101980
rect 197850 101910 198150 101980
rect 198350 101910 198650 101980
rect 198850 101910 199150 101980
rect 199350 101910 199650 101980
rect 199850 101910 200150 101980
rect 200350 101910 200650 101980
rect 200850 101910 201150 101980
rect 201350 101910 201650 101980
rect 201850 101910 202150 101980
rect 202350 101910 202650 101980
rect 202850 101910 203150 101980
rect 203350 101910 203650 101980
rect 203850 101910 204150 101980
rect 204350 101910 204650 101980
rect 204850 101910 205150 101980
rect 205350 101910 205650 101980
rect 205850 101910 206150 101980
rect 206350 101910 206650 101980
rect 206850 101910 207150 101980
rect 207350 101910 207650 101980
rect 207850 101910 208000 101980
rect 196000 101900 208000 101910
rect 196000 101880 196120 101900
rect 196380 101880 196620 101900
rect 196880 101880 197120 101900
rect 197380 101880 197620 101900
rect 197880 101880 198120 101900
rect 198380 101880 198620 101900
rect 198880 101880 199120 101900
rect 199380 101880 199620 101900
rect 199880 101880 200120 101900
rect 200380 101880 200620 101900
rect 200880 101880 201120 101900
rect 201380 101880 201620 101900
rect 201880 101880 202120 101900
rect 202380 101880 202620 101900
rect 202880 101880 203120 101900
rect 203380 101880 203620 101900
rect 203880 101880 204120 101900
rect 204380 101880 204620 101900
rect 204880 101880 205120 101900
rect 205380 101880 205620 101900
rect 205880 101880 206120 101900
rect 206380 101880 206620 101900
rect 206880 101880 207120 101900
rect 207380 101880 207620 101900
rect 207880 101880 208000 101900
rect 196000 101850 196100 101880
rect 196000 101650 196020 101850
rect 196090 101650 196100 101850
rect 196000 101620 196100 101650
rect 196400 101850 196600 101880
rect 196400 101650 196410 101850
rect 196480 101650 196520 101850
rect 196590 101650 196600 101850
rect 196400 101620 196600 101650
rect 196900 101850 197100 101880
rect 196900 101650 196910 101850
rect 196980 101650 197020 101850
rect 197090 101650 197100 101850
rect 196900 101620 197100 101650
rect 197400 101850 197600 101880
rect 197400 101650 197410 101850
rect 197480 101650 197520 101850
rect 197590 101650 197600 101850
rect 197400 101620 197600 101650
rect 197900 101850 198100 101880
rect 197900 101650 197910 101850
rect 197980 101650 198020 101850
rect 198090 101650 198100 101850
rect 197900 101620 198100 101650
rect 198400 101850 198600 101880
rect 198400 101650 198410 101850
rect 198480 101650 198520 101850
rect 198590 101650 198600 101850
rect 198400 101620 198600 101650
rect 198900 101850 199100 101880
rect 198900 101650 198910 101850
rect 198980 101650 199020 101850
rect 199090 101650 199100 101850
rect 198900 101620 199100 101650
rect 199400 101850 199600 101880
rect 199400 101650 199410 101850
rect 199480 101650 199520 101850
rect 199590 101650 199600 101850
rect 199400 101620 199600 101650
rect 199900 101850 200100 101880
rect 199900 101650 199910 101850
rect 199980 101650 200020 101850
rect 200090 101650 200100 101850
rect 199900 101620 200100 101650
rect 200400 101850 200600 101880
rect 200400 101650 200410 101850
rect 200480 101650 200520 101850
rect 200590 101650 200600 101850
rect 200400 101620 200600 101650
rect 200900 101850 201100 101880
rect 200900 101650 200910 101850
rect 200980 101650 201020 101850
rect 201090 101650 201100 101850
rect 200900 101620 201100 101650
rect 201400 101850 201600 101880
rect 201400 101650 201410 101850
rect 201480 101650 201520 101850
rect 201590 101650 201600 101850
rect 201400 101620 201600 101650
rect 201900 101850 202100 101880
rect 201900 101650 201910 101850
rect 201980 101650 202020 101850
rect 202090 101650 202100 101850
rect 201900 101620 202100 101650
rect 202400 101850 202600 101880
rect 202400 101650 202410 101850
rect 202480 101650 202520 101850
rect 202590 101650 202600 101850
rect 202400 101620 202600 101650
rect 202900 101850 203100 101880
rect 202900 101650 202910 101850
rect 202980 101650 203020 101850
rect 203090 101650 203100 101850
rect 202900 101620 203100 101650
rect 203400 101850 203600 101880
rect 203400 101650 203410 101850
rect 203480 101650 203520 101850
rect 203590 101650 203600 101850
rect 203400 101620 203600 101650
rect 203900 101850 204100 101880
rect 203900 101650 203910 101850
rect 203980 101650 204020 101850
rect 204090 101650 204100 101850
rect 203900 101620 204100 101650
rect 204400 101850 204600 101880
rect 204400 101650 204410 101850
rect 204480 101650 204520 101850
rect 204590 101650 204600 101850
rect 204400 101620 204600 101650
rect 204900 101850 205100 101880
rect 204900 101650 204910 101850
rect 204980 101650 205020 101850
rect 205090 101650 205100 101850
rect 204900 101620 205100 101650
rect 205400 101850 205600 101880
rect 205400 101650 205410 101850
rect 205480 101650 205520 101850
rect 205590 101650 205600 101850
rect 205400 101620 205600 101650
rect 205900 101850 206100 101880
rect 205900 101650 205910 101850
rect 205980 101650 206020 101850
rect 206090 101650 206100 101850
rect 205900 101620 206100 101650
rect 206400 101850 206600 101880
rect 206400 101650 206410 101850
rect 206480 101650 206520 101850
rect 206590 101650 206600 101850
rect 206400 101620 206600 101650
rect 206900 101850 207100 101880
rect 206900 101650 206910 101850
rect 206980 101650 207020 101850
rect 207090 101650 207100 101850
rect 206900 101620 207100 101650
rect 207400 101850 207600 101880
rect 207400 101650 207410 101850
rect 207480 101650 207520 101850
rect 207590 101650 207600 101850
rect 207400 101620 207600 101650
rect 207900 101850 208000 101880
rect 207900 101650 207910 101850
rect 207980 101650 208000 101850
rect 207900 101620 208000 101650
rect 196000 101600 196120 101620
rect 196380 101600 196620 101620
rect 196880 101600 197120 101620
rect 197380 101600 197620 101620
rect 197880 101600 198120 101620
rect 198380 101600 198620 101620
rect 198880 101600 199120 101620
rect 199380 101600 199620 101620
rect 199880 101600 200120 101620
rect 200380 101600 200620 101620
rect 200880 101600 201120 101620
rect 201380 101600 201620 101620
rect 201880 101600 202120 101620
rect 202380 101600 202620 101620
rect 202880 101600 203120 101620
rect 203380 101600 203620 101620
rect 203880 101600 204120 101620
rect 204380 101600 204620 101620
rect 204880 101600 205120 101620
rect 205380 101600 205620 101620
rect 205880 101600 206120 101620
rect 206380 101600 206620 101620
rect 206880 101600 207120 101620
rect 207380 101600 207620 101620
rect 207880 101600 208000 101620
rect 196000 101590 208000 101600
rect 196000 101520 196150 101590
rect 196350 101520 196650 101590
rect 196850 101520 197150 101590
rect 197350 101520 197650 101590
rect 197850 101520 198150 101590
rect 198350 101520 198650 101590
rect 198850 101520 199150 101590
rect 199350 101520 199650 101590
rect 199850 101520 200150 101590
rect 200350 101520 200650 101590
rect 200850 101520 201150 101590
rect 201350 101520 201650 101590
rect 201850 101520 202150 101590
rect 202350 101520 202650 101590
rect 202850 101520 203150 101590
rect 203350 101520 203650 101590
rect 203850 101520 204150 101590
rect 204350 101520 204650 101590
rect 204850 101520 205150 101590
rect 205350 101520 205650 101590
rect 205850 101520 206150 101590
rect 206350 101520 206650 101590
rect 206850 101520 207150 101590
rect 207350 101520 207650 101590
rect 207850 101520 208000 101590
rect 196000 101480 208000 101520
rect 196000 101410 196150 101480
rect 196350 101410 196650 101480
rect 196850 101410 197150 101480
rect 197350 101410 197650 101480
rect 197850 101410 198150 101480
rect 198350 101410 198650 101480
rect 198850 101410 199150 101480
rect 199350 101410 199650 101480
rect 199850 101410 200150 101480
rect 200350 101410 200650 101480
rect 200850 101410 201150 101480
rect 201350 101410 201650 101480
rect 201850 101410 202150 101480
rect 202350 101410 202650 101480
rect 202850 101410 203150 101480
rect 203350 101410 203650 101480
rect 203850 101410 204150 101480
rect 204350 101410 204650 101480
rect 204850 101410 205150 101480
rect 205350 101410 205650 101480
rect 205850 101410 206150 101480
rect 206350 101410 206650 101480
rect 206850 101410 207150 101480
rect 207350 101410 207650 101480
rect 207850 101410 208000 101480
rect 196000 101400 208000 101410
rect 196000 101380 196120 101400
rect 196380 101380 196620 101400
rect 196880 101380 197120 101400
rect 197380 101380 197620 101400
rect 197880 101380 198120 101400
rect 198380 101380 198620 101400
rect 198880 101380 199120 101400
rect 199380 101380 199620 101400
rect 199880 101380 200120 101400
rect 200380 101380 200620 101400
rect 200880 101380 201120 101400
rect 201380 101380 201620 101400
rect 201880 101380 202120 101400
rect 202380 101380 202620 101400
rect 202880 101380 203120 101400
rect 203380 101380 203620 101400
rect 203880 101380 204120 101400
rect 204380 101380 204620 101400
rect 204880 101380 205120 101400
rect 205380 101380 205620 101400
rect 205880 101380 206120 101400
rect 206380 101380 206620 101400
rect 206880 101380 207120 101400
rect 207380 101380 207620 101400
rect 207880 101380 208000 101400
rect 196000 101350 196100 101380
rect 196000 101150 196020 101350
rect 196090 101150 196100 101350
rect 196000 101120 196100 101150
rect 196400 101350 196600 101380
rect 196400 101150 196410 101350
rect 196480 101150 196520 101350
rect 196590 101150 196600 101350
rect 196400 101120 196600 101150
rect 196900 101350 197100 101380
rect 196900 101150 196910 101350
rect 196980 101150 197020 101350
rect 197090 101150 197100 101350
rect 196900 101120 197100 101150
rect 197400 101350 197600 101380
rect 197400 101150 197410 101350
rect 197480 101150 197520 101350
rect 197590 101150 197600 101350
rect 197400 101120 197600 101150
rect 197900 101350 198100 101380
rect 197900 101150 197910 101350
rect 197980 101150 198020 101350
rect 198090 101150 198100 101350
rect 197900 101120 198100 101150
rect 198400 101350 198600 101380
rect 198400 101150 198410 101350
rect 198480 101150 198520 101350
rect 198590 101150 198600 101350
rect 198400 101120 198600 101150
rect 198900 101350 199100 101380
rect 198900 101150 198910 101350
rect 198980 101150 199020 101350
rect 199090 101150 199100 101350
rect 198900 101120 199100 101150
rect 199400 101350 199600 101380
rect 199400 101150 199410 101350
rect 199480 101150 199520 101350
rect 199590 101150 199600 101350
rect 199400 101120 199600 101150
rect 199900 101350 200100 101380
rect 199900 101150 199910 101350
rect 199980 101150 200020 101350
rect 200090 101150 200100 101350
rect 199900 101120 200100 101150
rect 200400 101350 200600 101380
rect 200400 101150 200410 101350
rect 200480 101150 200520 101350
rect 200590 101150 200600 101350
rect 200400 101120 200600 101150
rect 200900 101350 201100 101380
rect 200900 101150 200910 101350
rect 200980 101150 201020 101350
rect 201090 101150 201100 101350
rect 200900 101120 201100 101150
rect 201400 101350 201600 101380
rect 201400 101150 201410 101350
rect 201480 101150 201520 101350
rect 201590 101150 201600 101350
rect 201400 101120 201600 101150
rect 201900 101350 202100 101380
rect 201900 101150 201910 101350
rect 201980 101150 202020 101350
rect 202090 101150 202100 101350
rect 201900 101120 202100 101150
rect 202400 101350 202600 101380
rect 202400 101150 202410 101350
rect 202480 101150 202520 101350
rect 202590 101150 202600 101350
rect 202400 101120 202600 101150
rect 202900 101350 203100 101380
rect 202900 101150 202910 101350
rect 202980 101150 203020 101350
rect 203090 101150 203100 101350
rect 202900 101120 203100 101150
rect 203400 101350 203600 101380
rect 203400 101150 203410 101350
rect 203480 101150 203520 101350
rect 203590 101150 203600 101350
rect 203400 101120 203600 101150
rect 203900 101350 204100 101380
rect 203900 101150 203910 101350
rect 203980 101150 204020 101350
rect 204090 101150 204100 101350
rect 203900 101120 204100 101150
rect 204400 101350 204600 101380
rect 204400 101150 204410 101350
rect 204480 101150 204520 101350
rect 204590 101150 204600 101350
rect 204400 101120 204600 101150
rect 204900 101350 205100 101380
rect 204900 101150 204910 101350
rect 204980 101150 205020 101350
rect 205090 101150 205100 101350
rect 204900 101120 205100 101150
rect 205400 101350 205600 101380
rect 205400 101150 205410 101350
rect 205480 101150 205520 101350
rect 205590 101150 205600 101350
rect 205400 101120 205600 101150
rect 205900 101350 206100 101380
rect 205900 101150 205910 101350
rect 205980 101150 206020 101350
rect 206090 101150 206100 101350
rect 205900 101120 206100 101150
rect 206400 101350 206600 101380
rect 206400 101150 206410 101350
rect 206480 101150 206520 101350
rect 206590 101150 206600 101350
rect 206400 101120 206600 101150
rect 206900 101350 207100 101380
rect 206900 101150 206910 101350
rect 206980 101150 207020 101350
rect 207090 101150 207100 101350
rect 206900 101120 207100 101150
rect 207400 101350 207600 101380
rect 207400 101150 207410 101350
rect 207480 101150 207520 101350
rect 207590 101150 207600 101350
rect 207400 101120 207600 101150
rect 207900 101350 208000 101380
rect 207900 101150 207910 101350
rect 207980 101150 208000 101350
rect 207900 101120 208000 101150
rect 196000 101100 196120 101120
rect 196380 101100 196620 101120
rect 196880 101100 197120 101120
rect 197380 101100 197620 101120
rect 197880 101100 198120 101120
rect 198380 101100 198620 101120
rect 198880 101100 199120 101120
rect 199380 101100 199620 101120
rect 199880 101100 200120 101120
rect 200380 101100 200620 101120
rect 200880 101100 201120 101120
rect 201380 101100 201620 101120
rect 201880 101100 202120 101120
rect 202380 101100 202620 101120
rect 202880 101100 203120 101120
rect 203380 101100 203620 101120
rect 203880 101100 204120 101120
rect 204380 101100 204620 101120
rect 204880 101100 205120 101120
rect 205380 101100 205620 101120
rect 205880 101100 206120 101120
rect 206380 101100 206620 101120
rect 206880 101100 207120 101120
rect 207380 101100 207620 101120
rect 207880 101100 208000 101120
rect 196000 101090 208000 101100
rect 196000 101020 196150 101090
rect 196350 101020 196650 101090
rect 196850 101020 197150 101090
rect 197350 101020 197650 101090
rect 197850 101020 198150 101090
rect 198350 101020 198650 101090
rect 198850 101020 199150 101090
rect 199350 101020 199650 101090
rect 199850 101020 200150 101090
rect 200350 101020 200650 101090
rect 200850 101020 201150 101090
rect 201350 101020 201650 101090
rect 201850 101020 202150 101090
rect 202350 101020 202650 101090
rect 202850 101020 203150 101090
rect 203350 101020 203650 101090
rect 203850 101020 204150 101090
rect 204350 101020 204650 101090
rect 204850 101020 205150 101090
rect 205350 101020 205650 101090
rect 205850 101020 206150 101090
rect 206350 101020 206650 101090
rect 206850 101020 207150 101090
rect 207350 101020 207650 101090
rect 207850 101020 208000 101090
rect 196000 100980 208000 101020
rect 196000 100910 196150 100980
rect 196350 100910 196650 100980
rect 196850 100910 197150 100980
rect 197350 100910 197650 100980
rect 197850 100910 198150 100980
rect 198350 100910 198650 100980
rect 198850 100910 199150 100980
rect 199350 100910 199650 100980
rect 199850 100910 200150 100980
rect 200350 100910 200650 100980
rect 200850 100910 201150 100980
rect 201350 100910 201650 100980
rect 201850 100910 202150 100980
rect 202350 100910 202650 100980
rect 202850 100910 203150 100980
rect 203350 100910 203650 100980
rect 203850 100910 204150 100980
rect 204350 100910 204650 100980
rect 204850 100910 205150 100980
rect 205350 100910 205650 100980
rect 205850 100910 206150 100980
rect 206350 100910 206650 100980
rect 206850 100910 207150 100980
rect 207350 100910 207650 100980
rect 207850 100910 208000 100980
rect 196000 100900 208000 100910
rect 196000 100880 196120 100900
rect 196380 100880 196620 100900
rect 196880 100880 197120 100900
rect 197380 100880 197620 100900
rect 197880 100880 198120 100900
rect 198380 100880 198620 100900
rect 198880 100880 199120 100900
rect 199380 100880 199620 100900
rect 199880 100880 200120 100900
rect 200380 100880 200620 100900
rect 200880 100880 201120 100900
rect 201380 100880 201620 100900
rect 201880 100880 202120 100900
rect 202380 100880 202620 100900
rect 202880 100880 203120 100900
rect 203380 100880 203620 100900
rect 203880 100880 204120 100900
rect 204380 100880 204620 100900
rect 204880 100880 205120 100900
rect 205380 100880 205620 100900
rect 205880 100880 206120 100900
rect 206380 100880 206620 100900
rect 206880 100880 207120 100900
rect 207380 100880 207620 100900
rect 207880 100880 208000 100900
rect 196000 100850 196100 100880
rect 196000 100650 196020 100850
rect 196090 100650 196100 100850
rect 196000 100620 196100 100650
rect 196400 100850 196600 100880
rect 196400 100650 196410 100850
rect 196480 100650 196520 100850
rect 196590 100650 196600 100850
rect 196400 100620 196600 100650
rect 196900 100850 197100 100880
rect 196900 100650 196910 100850
rect 196980 100650 197020 100850
rect 197090 100650 197100 100850
rect 196900 100620 197100 100650
rect 197400 100850 197600 100880
rect 197400 100650 197410 100850
rect 197480 100650 197520 100850
rect 197590 100650 197600 100850
rect 197400 100620 197600 100650
rect 197900 100850 198100 100880
rect 197900 100650 197910 100850
rect 197980 100650 198020 100850
rect 198090 100650 198100 100850
rect 197900 100620 198100 100650
rect 198400 100850 198600 100880
rect 198400 100650 198410 100850
rect 198480 100650 198520 100850
rect 198590 100650 198600 100850
rect 198400 100620 198600 100650
rect 198900 100850 199100 100880
rect 198900 100650 198910 100850
rect 198980 100650 199020 100850
rect 199090 100650 199100 100850
rect 198900 100620 199100 100650
rect 199400 100850 199600 100880
rect 199400 100650 199410 100850
rect 199480 100650 199520 100850
rect 199590 100650 199600 100850
rect 199400 100620 199600 100650
rect 199900 100850 200100 100880
rect 199900 100650 199910 100850
rect 199980 100650 200020 100850
rect 200090 100650 200100 100850
rect 199900 100620 200100 100650
rect 200400 100850 200600 100880
rect 200400 100650 200410 100850
rect 200480 100650 200520 100850
rect 200590 100650 200600 100850
rect 200400 100620 200600 100650
rect 200900 100850 201100 100880
rect 200900 100650 200910 100850
rect 200980 100650 201020 100850
rect 201090 100650 201100 100850
rect 200900 100620 201100 100650
rect 201400 100850 201600 100880
rect 201400 100650 201410 100850
rect 201480 100650 201520 100850
rect 201590 100650 201600 100850
rect 201400 100620 201600 100650
rect 201900 100850 202100 100880
rect 201900 100650 201910 100850
rect 201980 100650 202020 100850
rect 202090 100650 202100 100850
rect 201900 100620 202100 100650
rect 202400 100850 202600 100880
rect 202400 100650 202410 100850
rect 202480 100650 202520 100850
rect 202590 100650 202600 100850
rect 202400 100620 202600 100650
rect 202900 100850 203100 100880
rect 202900 100650 202910 100850
rect 202980 100650 203020 100850
rect 203090 100650 203100 100850
rect 202900 100620 203100 100650
rect 203400 100850 203600 100880
rect 203400 100650 203410 100850
rect 203480 100650 203520 100850
rect 203590 100650 203600 100850
rect 203400 100620 203600 100650
rect 203900 100850 204100 100880
rect 203900 100650 203910 100850
rect 203980 100650 204020 100850
rect 204090 100650 204100 100850
rect 203900 100620 204100 100650
rect 204400 100850 204600 100880
rect 204400 100650 204410 100850
rect 204480 100650 204520 100850
rect 204590 100650 204600 100850
rect 204400 100620 204600 100650
rect 204900 100850 205100 100880
rect 204900 100650 204910 100850
rect 204980 100650 205020 100850
rect 205090 100650 205100 100850
rect 204900 100620 205100 100650
rect 205400 100850 205600 100880
rect 205400 100650 205410 100850
rect 205480 100650 205520 100850
rect 205590 100650 205600 100850
rect 205400 100620 205600 100650
rect 205900 100850 206100 100880
rect 205900 100650 205910 100850
rect 205980 100650 206020 100850
rect 206090 100650 206100 100850
rect 205900 100620 206100 100650
rect 206400 100850 206600 100880
rect 206400 100650 206410 100850
rect 206480 100650 206520 100850
rect 206590 100650 206600 100850
rect 206400 100620 206600 100650
rect 206900 100850 207100 100880
rect 206900 100650 206910 100850
rect 206980 100650 207020 100850
rect 207090 100650 207100 100850
rect 206900 100620 207100 100650
rect 207400 100850 207600 100880
rect 207400 100650 207410 100850
rect 207480 100650 207520 100850
rect 207590 100650 207600 100850
rect 207400 100620 207600 100650
rect 207900 100850 208000 100880
rect 207900 100650 207910 100850
rect 207980 100650 208000 100850
rect 207900 100620 208000 100650
rect 196000 100600 196120 100620
rect 196380 100600 196620 100620
rect 196880 100600 197120 100620
rect 197380 100600 197620 100620
rect 197880 100600 198120 100620
rect 198380 100600 198620 100620
rect 198880 100600 199120 100620
rect 199380 100600 199620 100620
rect 199880 100600 200120 100620
rect 200380 100600 200620 100620
rect 200880 100600 201120 100620
rect 201380 100600 201620 100620
rect 201880 100600 202120 100620
rect 202380 100600 202620 100620
rect 202880 100600 203120 100620
rect 203380 100600 203620 100620
rect 203880 100600 204120 100620
rect 204380 100600 204620 100620
rect 204880 100600 205120 100620
rect 205380 100600 205620 100620
rect 205880 100600 206120 100620
rect 206380 100600 206620 100620
rect 206880 100600 207120 100620
rect 207380 100600 207620 100620
rect 207880 100600 208000 100620
rect 196000 100590 208000 100600
rect 196000 100520 196150 100590
rect 196350 100520 196650 100590
rect 196850 100520 197150 100590
rect 197350 100520 197650 100590
rect 197850 100520 198150 100590
rect 198350 100520 198650 100590
rect 198850 100520 199150 100590
rect 199350 100520 199650 100590
rect 199850 100520 200150 100590
rect 200350 100520 200650 100590
rect 200850 100520 201150 100590
rect 201350 100520 201650 100590
rect 201850 100520 202150 100590
rect 202350 100520 202650 100590
rect 202850 100520 203150 100590
rect 203350 100520 203650 100590
rect 203850 100520 204150 100590
rect 204350 100520 204650 100590
rect 204850 100520 205150 100590
rect 205350 100520 205650 100590
rect 205850 100520 206150 100590
rect 206350 100520 206650 100590
rect 206850 100520 207150 100590
rect 207350 100520 207650 100590
rect 207850 100520 208000 100590
rect 196000 100480 208000 100520
rect 196000 100410 196150 100480
rect 196350 100410 196650 100480
rect 196850 100410 197150 100480
rect 197350 100410 197650 100480
rect 197850 100410 198150 100480
rect 198350 100410 198650 100480
rect 198850 100410 199150 100480
rect 199350 100410 199650 100480
rect 199850 100410 200150 100480
rect 200350 100410 200650 100480
rect 200850 100410 201150 100480
rect 201350 100410 201650 100480
rect 201850 100410 202150 100480
rect 202350 100410 202650 100480
rect 202850 100410 203150 100480
rect 203350 100410 203650 100480
rect 203850 100410 204150 100480
rect 204350 100410 204650 100480
rect 204850 100410 205150 100480
rect 205350 100410 205650 100480
rect 205850 100410 206150 100480
rect 206350 100410 206650 100480
rect 206850 100410 207150 100480
rect 207350 100410 207650 100480
rect 207850 100410 208000 100480
rect 196000 100400 208000 100410
rect 196000 100380 196120 100400
rect 196380 100380 196620 100400
rect 196880 100380 197120 100400
rect 197380 100380 197620 100400
rect 197880 100380 198120 100400
rect 198380 100380 198620 100400
rect 198880 100380 199120 100400
rect 199380 100380 199620 100400
rect 199880 100380 200120 100400
rect 200380 100380 200620 100400
rect 200880 100380 201120 100400
rect 201380 100380 201620 100400
rect 201880 100380 202120 100400
rect 202380 100380 202620 100400
rect 202880 100380 203120 100400
rect 203380 100380 203620 100400
rect 203880 100380 204120 100400
rect 204380 100380 204620 100400
rect 204880 100380 205120 100400
rect 205380 100380 205620 100400
rect 205880 100380 206120 100400
rect 206380 100380 206620 100400
rect 206880 100380 207120 100400
rect 207380 100380 207620 100400
rect 207880 100380 208000 100400
rect 196000 100350 196100 100380
rect 196000 100150 196020 100350
rect 196090 100150 196100 100350
rect 196000 100120 196100 100150
rect 196400 100350 196600 100380
rect 196400 100150 196410 100350
rect 196480 100150 196520 100350
rect 196590 100150 196600 100350
rect 196400 100120 196600 100150
rect 196900 100350 197100 100380
rect 196900 100150 196910 100350
rect 196980 100150 197020 100350
rect 197090 100150 197100 100350
rect 196900 100120 197100 100150
rect 197400 100350 197600 100380
rect 197400 100150 197410 100350
rect 197480 100150 197520 100350
rect 197590 100150 197600 100350
rect 197400 100120 197600 100150
rect 197900 100350 198100 100380
rect 197900 100150 197910 100350
rect 197980 100150 198020 100350
rect 198090 100150 198100 100350
rect 197900 100120 198100 100150
rect 198400 100350 198600 100380
rect 198400 100150 198410 100350
rect 198480 100150 198520 100350
rect 198590 100150 198600 100350
rect 198400 100120 198600 100150
rect 198900 100350 199100 100380
rect 198900 100150 198910 100350
rect 198980 100150 199020 100350
rect 199090 100150 199100 100350
rect 198900 100120 199100 100150
rect 199400 100350 199600 100380
rect 199400 100150 199410 100350
rect 199480 100150 199520 100350
rect 199590 100150 199600 100350
rect 199400 100120 199600 100150
rect 199900 100350 200100 100380
rect 199900 100150 199910 100350
rect 199980 100150 200020 100350
rect 200090 100150 200100 100350
rect 199900 100120 200100 100150
rect 200400 100350 200600 100380
rect 200400 100150 200410 100350
rect 200480 100150 200520 100350
rect 200590 100150 200600 100350
rect 200400 100120 200600 100150
rect 200900 100350 201100 100380
rect 200900 100150 200910 100350
rect 200980 100150 201020 100350
rect 201090 100150 201100 100350
rect 200900 100120 201100 100150
rect 201400 100350 201600 100380
rect 201400 100150 201410 100350
rect 201480 100150 201520 100350
rect 201590 100150 201600 100350
rect 201400 100120 201600 100150
rect 201900 100350 202100 100380
rect 201900 100150 201910 100350
rect 201980 100150 202020 100350
rect 202090 100150 202100 100350
rect 201900 100120 202100 100150
rect 202400 100350 202600 100380
rect 202400 100150 202410 100350
rect 202480 100150 202520 100350
rect 202590 100150 202600 100350
rect 202400 100120 202600 100150
rect 202900 100350 203100 100380
rect 202900 100150 202910 100350
rect 202980 100150 203020 100350
rect 203090 100150 203100 100350
rect 202900 100120 203100 100150
rect 203400 100350 203600 100380
rect 203400 100150 203410 100350
rect 203480 100150 203520 100350
rect 203590 100150 203600 100350
rect 203400 100120 203600 100150
rect 203900 100350 204100 100380
rect 203900 100150 203910 100350
rect 203980 100150 204020 100350
rect 204090 100150 204100 100350
rect 203900 100120 204100 100150
rect 204400 100350 204600 100380
rect 204400 100150 204410 100350
rect 204480 100150 204520 100350
rect 204590 100150 204600 100350
rect 204400 100120 204600 100150
rect 204900 100350 205100 100380
rect 204900 100150 204910 100350
rect 204980 100150 205020 100350
rect 205090 100150 205100 100350
rect 204900 100120 205100 100150
rect 205400 100350 205600 100380
rect 205400 100150 205410 100350
rect 205480 100150 205520 100350
rect 205590 100150 205600 100350
rect 205400 100120 205600 100150
rect 205900 100350 206100 100380
rect 205900 100150 205910 100350
rect 205980 100150 206020 100350
rect 206090 100150 206100 100350
rect 205900 100120 206100 100150
rect 206400 100350 206600 100380
rect 206400 100150 206410 100350
rect 206480 100150 206520 100350
rect 206590 100150 206600 100350
rect 206400 100120 206600 100150
rect 206900 100350 207100 100380
rect 206900 100150 206910 100350
rect 206980 100150 207020 100350
rect 207090 100150 207100 100350
rect 206900 100120 207100 100150
rect 207400 100350 207600 100380
rect 207400 100150 207410 100350
rect 207480 100150 207520 100350
rect 207590 100150 207600 100350
rect 207400 100120 207600 100150
rect 207900 100350 208000 100380
rect 207900 100150 207910 100350
rect 207980 100150 208000 100350
rect 207900 100120 208000 100150
rect 196000 100100 196120 100120
rect 196380 100100 196620 100120
rect 196880 100100 197120 100120
rect 197380 100100 197620 100120
rect 197880 100100 198120 100120
rect 198380 100100 198620 100120
rect 198880 100100 199120 100120
rect 199380 100100 199620 100120
rect 199880 100100 200120 100120
rect 200380 100100 200620 100120
rect 200880 100100 201120 100120
rect 201380 100100 201620 100120
rect 201880 100100 202120 100120
rect 202380 100100 202620 100120
rect 202880 100100 203120 100120
rect 203380 100100 203620 100120
rect 203880 100100 204120 100120
rect 204380 100100 204620 100120
rect 204880 100100 205120 100120
rect 205380 100100 205620 100120
rect 205880 100100 206120 100120
rect 206380 100100 206620 100120
rect 206880 100100 207120 100120
rect 207380 100100 207620 100120
rect 207880 100100 208000 100120
rect 196000 100090 208000 100100
rect 196000 100020 196150 100090
rect 196350 100020 196650 100090
rect 196850 100020 197150 100090
rect 197350 100020 197650 100090
rect 197850 100020 198150 100090
rect 198350 100020 198650 100090
rect 198850 100020 199150 100090
rect 199350 100020 199650 100090
rect 199850 100020 200150 100090
rect 200350 100020 200650 100090
rect 200850 100020 201150 100090
rect 201350 100020 201650 100090
rect 201850 100020 202150 100090
rect 202350 100020 202650 100090
rect 202850 100020 203150 100090
rect 203350 100020 203650 100090
rect 203850 100020 204150 100090
rect 204350 100020 204650 100090
rect 204850 100020 205150 100090
rect 205350 100020 205650 100090
rect 205850 100020 206150 100090
rect 206350 100020 206650 100090
rect 206850 100020 207150 100090
rect 207350 100020 207650 100090
rect 207850 100020 208000 100090
rect 196000 99980 208000 100020
rect 196000 99910 196150 99980
rect 196350 99910 196650 99980
rect 196850 99910 197150 99980
rect 197350 99910 197650 99980
rect 197850 99910 198150 99980
rect 198350 99910 198650 99980
rect 198850 99910 199150 99980
rect 199350 99910 199650 99980
rect 199850 99910 200150 99980
rect 200350 99910 200650 99980
rect 200850 99910 201150 99980
rect 201350 99910 201650 99980
rect 201850 99910 202150 99980
rect 202350 99910 202650 99980
rect 202850 99910 203150 99980
rect 203350 99910 203650 99980
rect 203850 99910 204150 99980
rect 204350 99910 204650 99980
rect 204850 99910 205150 99980
rect 205350 99910 205650 99980
rect 205850 99910 206150 99980
rect 206350 99910 206650 99980
rect 206850 99910 207150 99980
rect 207350 99910 207650 99980
rect 207850 99910 208000 99980
rect 196000 99900 208000 99910
rect 196000 99880 196120 99900
rect 196380 99880 196620 99900
rect 196880 99880 197120 99900
rect 197380 99880 197620 99900
rect 197880 99880 198120 99900
rect 198380 99880 198620 99900
rect 198880 99880 199120 99900
rect 199380 99880 199620 99900
rect 199880 99880 200120 99900
rect 200380 99880 200620 99900
rect 200880 99880 201120 99900
rect 201380 99880 201620 99900
rect 201880 99880 202120 99900
rect 202380 99880 202620 99900
rect 202880 99880 203120 99900
rect 203380 99880 203620 99900
rect 203880 99880 204120 99900
rect 204380 99880 204620 99900
rect 204880 99880 205120 99900
rect 205380 99880 205620 99900
rect 205880 99880 206120 99900
rect 206380 99880 206620 99900
rect 206880 99880 207120 99900
rect 207380 99880 207620 99900
rect 207880 99880 208000 99900
rect 196000 99850 196100 99880
rect 196000 99650 196020 99850
rect 196090 99650 196100 99850
rect 196000 99620 196100 99650
rect 196400 99850 196600 99880
rect 196400 99650 196410 99850
rect 196480 99650 196520 99850
rect 196590 99650 196600 99850
rect 196400 99620 196600 99650
rect 196900 99850 197100 99880
rect 196900 99650 196910 99850
rect 196980 99650 197020 99850
rect 197090 99650 197100 99850
rect 196900 99620 197100 99650
rect 197400 99850 197600 99880
rect 197400 99650 197410 99850
rect 197480 99650 197520 99850
rect 197590 99650 197600 99850
rect 197400 99620 197600 99650
rect 197900 99850 198100 99880
rect 197900 99650 197910 99850
rect 197980 99650 198020 99850
rect 198090 99650 198100 99850
rect 197900 99620 198100 99650
rect 198400 99850 198600 99880
rect 198400 99650 198410 99850
rect 198480 99650 198520 99850
rect 198590 99650 198600 99850
rect 198400 99620 198600 99650
rect 198900 99850 199100 99880
rect 198900 99650 198910 99850
rect 198980 99650 199020 99850
rect 199090 99650 199100 99850
rect 198900 99620 199100 99650
rect 199400 99850 199600 99880
rect 199400 99650 199410 99850
rect 199480 99650 199520 99850
rect 199590 99650 199600 99850
rect 199400 99620 199600 99650
rect 199900 99850 200100 99880
rect 199900 99650 199910 99850
rect 199980 99650 200020 99850
rect 200090 99650 200100 99850
rect 199900 99620 200100 99650
rect 200400 99850 200600 99880
rect 200400 99650 200410 99850
rect 200480 99650 200520 99850
rect 200590 99650 200600 99850
rect 200400 99620 200600 99650
rect 200900 99850 201100 99880
rect 200900 99650 200910 99850
rect 200980 99650 201020 99850
rect 201090 99650 201100 99850
rect 200900 99620 201100 99650
rect 201400 99850 201600 99880
rect 201400 99650 201410 99850
rect 201480 99650 201520 99850
rect 201590 99650 201600 99850
rect 201400 99620 201600 99650
rect 201900 99850 202100 99880
rect 201900 99650 201910 99850
rect 201980 99650 202020 99850
rect 202090 99650 202100 99850
rect 201900 99620 202100 99650
rect 202400 99850 202600 99880
rect 202400 99650 202410 99850
rect 202480 99650 202520 99850
rect 202590 99650 202600 99850
rect 202400 99620 202600 99650
rect 202900 99850 203100 99880
rect 202900 99650 202910 99850
rect 202980 99650 203020 99850
rect 203090 99650 203100 99850
rect 202900 99620 203100 99650
rect 203400 99850 203600 99880
rect 203400 99650 203410 99850
rect 203480 99650 203520 99850
rect 203590 99650 203600 99850
rect 203400 99620 203600 99650
rect 203900 99850 204100 99880
rect 203900 99650 203910 99850
rect 203980 99650 204020 99850
rect 204090 99650 204100 99850
rect 203900 99620 204100 99650
rect 204400 99850 204600 99880
rect 204400 99650 204410 99850
rect 204480 99650 204520 99850
rect 204590 99650 204600 99850
rect 204400 99620 204600 99650
rect 204900 99850 205100 99880
rect 204900 99650 204910 99850
rect 204980 99650 205020 99850
rect 205090 99650 205100 99850
rect 204900 99620 205100 99650
rect 205400 99850 205600 99880
rect 205400 99650 205410 99850
rect 205480 99650 205520 99850
rect 205590 99650 205600 99850
rect 205400 99620 205600 99650
rect 205900 99850 206100 99880
rect 205900 99650 205910 99850
rect 205980 99650 206020 99850
rect 206090 99650 206100 99850
rect 205900 99620 206100 99650
rect 206400 99850 206600 99880
rect 206400 99650 206410 99850
rect 206480 99650 206520 99850
rect 206590 99650 206600 99850
rect 206400 99620 206600 99650
rect 206900 99850 207100 99880
rect 206900 99650 206910 99850
rect 206980 99650 207020 99850
rect 207090 99650 207100 99850
rect 206900 99620 207100 99650
rect 207400 99850 207600 99880
rect 207400 99650 207410 99850
rect 207480 99650 207520 99850
rect 207590 99650 207600 99850
rect 207400 99620 207600 99650
rect 207900 99850 208000 99880
rect 207900 99650 207910 99850
rect 207980 99650 208000 99850
rect 207900 99620 208000 99650
rect 196000 99600 196120 99620
rect 196380 99600 196620 99620
rect 196880 99600 197120 99620
rect 197380 99600 197620 99620
rect 197880 99600 198120 99620
rect 198380 99600 198620 99620
rect 198880 99600 199120 99620
rect 199380 99600 199620 99620
rect 199880 99600 200120 99620
rect 200380 99600 200620 99620
rect 200880 99600 201120 99620
rect 201380 99600 201620 99620
rect 201880 99600 202120 99620
rect 202380 99600 202620 99620
rect 202880 99600 203120 99620
rect 203380 99600 203620 99620
rect 203880 99600 204120 99620
rect 204380 99600 204620 99620
rect 204880 99600 205120 99620
rect 205380 99600 205620 99620
rect 205880 99600 206120 99620
rect 206380 99600 206620 99620
rect 206880 99600 207120 99620
rect 207380 99600 207620 99620
rect 207880 99600 208000 99620
rect 196000 99590 208000 99600
rect 196000 99520 196150 99590
rect 196350 99520 196650 99590
rect 196850 99520 197150 99590
rect 197350 99520 197650 99590
rect 197850 99520 198150 99590
rect 198350 99520 198650 99590
rect 198850 99520 199150 99590
rect 199350 99520 199650 99590
rect 199850 99520 200150 99590
rect 200350 99520 200650 99590
rect 200850 99520 201150 99590
rect 201350 99520 201650 99590
rect 201850 99520 202150 99590
rect 202350 99520 202650 99590
rect 202850 99520 203150 99590
rect 203350 99520 203650 99590
rect 203850 99520 204150 99590
rect 204350 99520 204650 99590
rect 204850 99520 205150 99590
rect 205350 99520 205650 99590
rect 205850 99520 206150 99590
rect 206350 99520 206650 99590
rect 206850 99520 207150 99590
rect 207350 99520 207650 99590
rect 207850 99520 208000 99590
rect 196000 99480 208000 99520
rect 196000 99410 196150 99480
rect 196350 99410 196650 99480
rect 196850 99410 197150 99480
rect 197350 99410 197650 99480
rect 197850 99410 198150 99480
rect 198350 99410 198650 99480
rect 198850 99410 199150 99480
rect 199350 99410 199650 99480
rect 199850 99410 200150 99480
rect 200350 99410 200650 99480
rect 200850 99410 201150 99480
rect 201350 99410 201650 99480
rect 201850 99410 202150 99480
rect 202350 99410 202650 99480
rect 202850 99410 203150 99480
rect 203350 99410 203650 99480
rect 203850 99410 204150 99480
rect 204350 99410 204650 99480
rect 204850 99410 205150 99480
rect 205350 99410 205650 99480
rect 205850 99410 206150 99480
rect 206350 99410 206650 99480
rect 206850 99410 207150 99480
rect 207350 99410 207650 99480
rect 207850 99410 208000 99480
rect 196000 99400 208000 99410
rect 196000 99380 196120 99400
rect 196380 99380 196620 99400
rect 196880 99380 197120 99400
rect 197380 99380 197620 99400
rect 197880 99380 198120 99400
rect 198380 99380 198620 99400
rect 198880 99380 199120 99400
rect 199380 99380 199620 99400
rect 199880 99380 200120 99400
rect 200380 99380 200620 99400
rect 200880 99380 201120 99400
rect 201380 99380 201620 99400
rect 201880 99380 202120 99400
rect 202380 99380 202620 99400
rect 202880 99380 203120 99400
rect 203380 99380 203620 99400
rect 203880 99380 204120 99400
rect 204380 99380 204620 99400
rect 204880 99380 205120 99400
rect 205380 99380 205620 99400
rect 205880 99380 206120 99400
rect 206380 99380 206620 99400
rect 206880 99380 207120 99400
rect 207380 99380 207620 99400
rect 207880 99380 208000 99400
rect 196000 99350 196100 99380
rect 196000 99150 196020 99350
rect 196090 99150 196100 99350
rect 196000 99120 196100 99150
rect 196400 99350 196600 99380
rect 196400 99150 196410 99350
rect 196480 99150 196520 99350
rect 196590 99150 196600 99350
rect 196400 99120 196600 99150
rect 196900 99350 197100 99380
rect 196900 99150 196910 99350
rect 196980 99150 197020 99350
rect 197090 99150 197100 99350
rect 196900 99120 197100 99150
rect 197400 99350 197600 99380
rect 197400 99150 197410 99350
rect 197480 99150 197520 99350
rect 197590 99150 197600 99350
rect 197400 99120 197600 99150
rect 197900 99350 198100 99380
rect 197900 99150 197910 99350
rect 197980 99150 198020 99350
rect 198090 99150 198100 99350
rect 197900 99120 198100 99150
rect 198400 99350 198600 99380
rect 198400 99150 198410 99350
rect 198480 99150 198520 99350
rect 198590 99150 198600 99350
rect 198400 99120 198600 99150
rect 198900 99350 199100 99380
rect 198900 99150 198910 99350
rect 198980 99150 199020 99350
rect 199090 99150 199100 99350
rect 198900 99120 199100 99150
rect 199400 99350 199600 99380
rect 199400 99150 199410 99350
rect 199480 99150 199520 99350
rect 199590 99150 199600 99350
rect 199400 99120 199600 99150
rect 199900 99350 200100 99380
rect 199900 99150 199910 99350
rect 199980 99150 200020 99350
rect 200090 99150 200100 99350
rect 199900 99120 200100 99150
rect 200400 99350 200600 99380
rect 200400 99150 200410 99350
rect 200480 99150 200520 99350
rect 200590 99150 200600 99350
rect 200400 99120 200600 99150
rect 200900 99350 201100 99380
rect 200900 99150 200910 99350
rect 200980 99150 201020 99350
rect 201090 99150 201100 99350
rect 200900 99120 201100 99150
rect 201400 99350 201600 99380
rect 201400 99150 201410 99350
rect 201480 99150 201520 99350
rect 201590 99150 201600 99350
rect 201400 99120 201600 99150
rect 201900 99350 202100 99380
rect 201900 99150 201910 99350
rect 201980 99150 202020 99350
rect 202090 99150 202100 99350
rect 201900 99120 202100 99150
rect 202400 99350 202600 99380
rect 202400 99150 202410 99350
rect 202480 99150 202520 99350
rect 202590 99150 202600 99350
rect 202400 99120 202600 99150
rect 202900 99350 203100 99380
rect 202900 99150 202910 99350
rect 202980 99150 203020 99350
rect 203090 99150 203100 99350
rect 202900 99120 203100 99150
rect 203400 99350 203600 99380
rect 203400 99150 203410 99350
rect 203480 99150 203520 99350
rect 203590 99150 203600 99350
rect 203400 99120 203600 99150
rect 203900 99350 204100 99380
rect 203900 99150 203910 99350
rect 203980 99150 204020 99350
rect 204090 99150 204100 99350
rect 203900 99120 204100 99150
rect 204400 99350 204600 99380
rect 204400 99150 204410 99350
rect 204480 99150 204520 99350
rect 204590 99150 204600 99350
rect 204400 99120 204600 99150
rect 204900 99350 205100 99380
rect 204900 99150 204910 99350
rect 204980 99150 205020 99350
rect 205090 99150 205100 99350
rect 204900 99120 205100 99150
rect 205400 99350 205600 99380
rect 205400 99150 205410 99350
rect 205480 99150 205520 99350
rect 205590 99150 205600 99350
rect 205400 99120 205600 99150
rect 205900 99350 206100 99380
rect 205900 99150 205910 99350
rect 205980 99150 206020 99350
rect 206090 99150 206100 99350
rect 205900 99120 206100 99150
rect 206400 99350 206600 99380
rect 206400 99150 206410 99350
rect 206480 99150 206520 99350
rect 206590 99150 206600 99350
rect 206400 99120 206600 99150
rect 206900 99350 207100 99380
rect 206900 99150 206910 99350
rect 206980 99150 207020 99350
rect 207090 99150 207100 99350
rect 206900 99120 207100 99150
rect 207400 99350 207600 99380
rect 207400 99150 207410 99350
rect 207480 99150 207520 99350
rect 207590 99150 207600 99350
rect 207400 99120 207600 99150
rect 207900 99350 208000 99380
rect 207900 99150 207910 99350
rect 207980 99150 208000 99350
rect 207900 99120 208000 99150
rect 196000 99100 196120 99120
rect 196380 99100 196620 99120
rect 196880 99100 197120 99120
rect 197380 99100 197620 99120
rect 197880 99100 198120 99120
rect 198380 99100 198620 99120
rect 198880 99100 199120 99120
rect 199380 99100 199620 99120
rect 199880 99100 200120 99120
rect 200380 99100 200620 99120
rect 200880 99100 201120 99120
rect 201380 99100 201620 99120
rect 201880 99100 202120 99120
rect 202380 99100 202620 99120
rect 202880 99100 203120 99120
rect 203380 99100 203620 99120
rect 203880 99100 204120 99120
rect 204380 99100 204620 99120
rect 204880 99100 205120 99120
rect 205380 99100 205620 99120
rect 205880 99100 206120 99120
rect 206380 99100 206620 99120
rect 206880 99100 207120 99120
rect 207380 99100 207620 99120
rect 207880 99100 208000 99120
rect 196000 99090 208000 99100
rect 196000 99020 196150 99090
rect 196350 99020 196650 99090
rect 196850 99020 197150 99090
rect 197350 99020 197650 99090
rect 197850 99020 198150 99090
rect 198350 99020 198650 99090
rect 198850 99020 199150 99090
rect 199350 99020 199650 99090
rect 199850 99020 200150 99090
rect 200350 99020 200650 99090
rect 200850 99020 201150 99090
rect 201350 99020 201650 99090
rect 201850 99020 202150 99090
rect 202350 99020 202650 99090
rect 202850 99020 203150 99090
rect 203350 99020 203650 99090
rect 203850 99020 204150 99090
rect 204350 99020 204650 99090
rect 204850 99020 205150 99090
rect 205350 99020 205650 99090
rect 205850 99020 206150 99090
rect 206350 99020 206650 99090
rect 206850 99020 207150 99090
rect 207350 99020 207650 99090
rect 207850 99020 208000 99090
rect 196000 98980 208000 99020
rect 196000 98910 196150 98980
rect 196350 98910 196650 98980
rect 196850 98910 197150 98980
rect 197350 98910 197650 98980
rect 197850 98910 198150 98980
rect 198350 98910 198650 98980
rect 198850 98910 199150 98980
rect 199350 98910 199650 98980
rect 199850 98910 200150 98980
rect 200350 98910 200650 98980
rect 200850 98910 201150 98980
rect 201350 98910 201650 98980
rect 201850 98910 202150 98980
rect 202350 98910 202650 98980
rect 202850 98910 203150 98980
rect 203350 98910 203650 98980
rect 203850 98910 204150 98980
rect 204350 98910 204650 98980
rect 204850 98910 205150 98980
rect 205350 98910 205650 98980
rect 205850 98910 206150 98980
rect 206350 98910 206650 98980
rect 206850 98910 207150 98980
rect 207350 98910 207650 98980
rect 207850 98910 208000 98980
rect 196000 98900 208000 98910
rect 196000 98880 196120 98900
rect 196380 98880 196620 98900
rect 196880 98880 197120 98900
rect 197380 98880 197620 98900
rect 197880 98880 198120 98900
rect 198380 98880 198620 98900
rect 198880 98880 199120 98900
rect 199380 98880 199620 98900
rect 199880 98880 200120 98900
rect 200380 98880 200620 98900
rect 200880 98880 201120 98900
rect 201380 98880 201620 98900
rect 201880 98880 202120 98900
rect 202380 98880 202620 98900
rect 202880 98880 203120 98900
rect 203380 98880 203620 98900
rect 203880 98880 204120 98900
rect 204380 98880 204620 98900
rect 204880 98880 205120 98900
rect 205380 98880 205620 98900
rect 205880 98880 206120 98900
rect 206380 98880 206620 98900
rect 206880 98880 207120 98900
rect 207380 98880 207620 98900
rect 207880 98880 208000 98900
rect 196000 98850 196100 98880
rect 196000 98650 196020 98850
rect 196090 98650 196100 98850
rect 196000 98620 196100 98650
rect 196400 98850 196600 98880
rect 196400 98650 196410 98850
rect 196480 98650 196520 98850
rect 196590 98650 196600 98850
rect 196400 98620 196600 98650
rect 196900 98850 197100 98880
rect 196900 98650 196910 98850
rect 196980 98650 197020 98850
rect 197090 98650 197100 98850
rect 196900 98620 197100 98650
rect 197400 98850 197600 98880
rect 197400 98650 197410 98850
rect 197480 98650 197520 98850
rect 197590 98650 197600 98850
rect 197400 98620 197600 98650
rect 197900 98850 198100 98880
rect 197900 98650 197910 98850
rect 197980 98650 198020 98850
rect 198090 98650 198100 98850
rect 197900 98620 198100 98650
rect 198400 98850 198600 98880
rect 198400 98650 198410 98850
rect 198480 98650 198520 98850
rect 198590 98650 198600 98850
rect 198400 98620 198600 98650
rect 198900 98850 199100 98880
rect 198900 98650 198910 98850
rect 198980 98650 199020 98850
rect 199090 98650 199100 98850
rect 198900 98620 199100 98650
rect 199400 98850 199600 98880
rect 199400 98650 199410 98850
rect 199480 98650 199520 98850
rect 199590 98650 199600 98850
rect 199400 98620 199600 98650
rect 199900 98850 200100 98880
rect 199900 98650 199910 98850
rect 199980 98650 200020 98850
rect 200090 98650 200100 98850
rect 199900 98620 200100 98650
rect 200400 98850 200600 98880
rect 200400 98650 200410 98850
rect 200480 98650 200520 98850
rect 200590 98650 200600 98850
rect 200400 98620 200600 98650
rect 200900 98850 201100 98880
rect 200900 98650 200910 98850
rect 200980 98650 201020 98850
rect 201090 98650 201100 98850
rect 200900 98620 201100 98650
rect 201400 98850 201600 98880
rect 201400 98650 201410 98850
rect 201480 98650 201520 98850
rect 201590 98650 201600 98850
rect 201400 98620 201600 98650
rect 201900 98850 202100 98880
rect 201900 98650 201910 98850
rect 201980 98650 202020 98850
rect 202090 98650 202100 98850
rect 201900 98620 202100 98650
rect 202400 98850 202600 98880
rect 202400 98650 202410 98850
rect 202480 98650 202520 98850
rect 202590 98650 202600 98850
rect 202400 98620 202600 98650
rect 202900 98850 203100 98880
rect 202900 98650 202910 98850
rect 202980 98650 203020 98850
rect 203090 98650 203100 98850
rect 202900 98620 203100 98650
rect 203400 98850 203600 98880
rect 203400 98650 203410 98850
rect 203480 98650 203520 98850
rect 203590 98650 203600 98850
rect 203400 98620 203600 98650
rect 203900 98850 204100 98880
rect 203900 98650 203910 98850
rect 203980 98650 204020 98850
rect 204090 98650 204100 98850
rect 203900 98620 204100 98650
rect 204400 98850 204600 98880
rect 204400 98650 204410 98850
rect 204480 98650 204520 98850
rect 204590 98650 204600 98850
rect 204400 98620 204600 98650
rect 204900 98850 205100 98880
rect 204900 98650 204910 98850
rect 204980 98650 205020 98850
rect 205090 98650 205100 98850
rect 204900 98620 205100 98650
rect 205400 98850 205600 98880
rect 205400 98650 205410 98850
rect 205480 98650 205520 98850
rect 205590 98650 205600 98850
rect 205400 98620 205600 98650
rect 205900 98850 206100 98880
rect 205900 98650 205910 98850
rect 205980 98650 206020 98850
rect 206090 98650 206100 98850
rect 205900 98620 206100 98650
rect 206400 98850 206600 98880
rect 206400 98650 206410 98850
rect 206480 98650 206520 98850
rect 206590 98650 206600 98850
rect 206400 98620 206600 98650
rect 206900 98850 207100 98880
rect 206900 98650 206910 98850
rect 206980 98650 207020 98850
rect 207090 98650 207100 98850
rect 206900 98620 207100 98650
rect 207400 98850 207600 98880
rect 207400 98650 207410 98850
rect 207480 98650 207520 98850
rect 207590 98650 207600 98850
rect 207400 98620 207600 98650
rect 207900 98850 208000 98880
rect 207900 98650 207910 98850
rect 207980 98650 208000 98850
rect 207900 98620 208000 98650
rect 196000 98600 196120 98620
rect 196380 98600 196620 98620
rect 196880 98600 197120 98620
rect 197380 98600 197620 98620
rect 197880 98600 198120 98620
rect 198380 98600 198620 98620
rect 198880 98600 199120 98620
rect 199380 98600 199620 98620
rect 199880 98600 200120 98620
rect 200380 98600 200620 98620
rect 200880 98600 201120 98620
rect 201380 98600 201620 98620
rect 201880 98600 202120 98620
rect 202380 98600 202620 98620
rect 202880 98600 203120 98620
rect 203380 98600 203620 98620
rect 203880 98600 204120 98620
rect 204380 98600 204620 98620
rect 204880 98600 205120 98620
rect 205380 98600 205620 98620
rect 205880 98600 206120 98620
rect 206380 98600 206620 98620
rect 206880 98600 207120 98620
rect 207380 98600 207620 98620
rect 207880 98600 208000 98620
rect 196000 98590 208000 98600
rect 196000 98520 196150 98590
rect 196350 98520 196650 98590
rect 196850 98520 197150 98590
rect 197350 98520 197650 98590
rect 197850 98520 198150 98590
rect 198350 98520 198650 98590
rect 198850 98520 199150 98590
rect 199350 98520 199650 98590
rect 199850 98520 200150 98590
rect 200350 98520 200650 98590
rect 200850 98520 201150 98590
rect 201350 98520 201650 98590
rect 201850 98520 202150 98590
rect 202350 98520 202650 98590
rect 202850 98520 203150 98590
rect 203350 98520 203650 98590
rect 203850 98520 204150 98590
rect 204350 98520 204650 98590
rect 204850 98520 205150 98590
rect 205350 98520 205650 98590
rect 205850 98520 206150 98590
rect 206350 98520 206650 98590
rect 206850 98520 207150 98590
rect 207350 98520 207650 98590
rect 207850 98520 208000 98590
rect 196000 98480 208000 98520
rect 196000 98410 196150 98480
rect 196350 98410 196650 98480
rect 196850 98410 197150 98480
rect 197350 98410 197650 98480
rect 197850 98410 198150 98480
rect 198350 98410 198650 98480
rect 198850 98410 199150 98480
rect 199350 98410 199650 98480
rect 199850 98410 200150 98480
rect 200350 98410 200650 98480
rect 200850 98410 201150 98480
rect 201350 98410 201650 98480
rect 201850 98410 202150 98480
rect 202350 98410 202650 98480
rect 202850 98410 203150 98480
rect 203350 98410 203650 98480
rect 203850 98410 204150 98480
rect 204350 98410 204650 98480
rect 204850 98410 205150 98480
rect 205350 98410 205650 98480
rect 205850 98410 206150 98480
rect 206350 98410 206650 98480
rect 206850 98410 207150 98480
rect 207350 98410 207650 98480
rect 207850 98410 208000 98480
rect 196000 98400 208000 98410
rect 196000 98380 196120 98400
rect 196380 98380 196620 98400
rect 196880 98380 197120 98400
rect 197380 98380 197620 98400
rect 197880 98380 198120 98400
rect 198380 98380 198620 98400
rect 198880 98380 199120 98400
rect 199380 98380 199620 98400
rect 199880 98380 200120 98400
rect 200380 98380 200620 98400
rect 200880 98380 201120 98400
rect 201380 98380 201620 98400
rect 201880 98380 202120 98400
rect 202380 98380 202620 98400
rect 202880 98380 203120 98400
rect 203380 98380 203620 98400
rect 203880 98380 204120 98400
rect 204380 98380 204620 98400
rect 204880 98380 205120 98400
rect 205380 98380 205620 98400
rect 205880 98380 206120 98400
rect 206380 98380 206620 98400
rect 206880 98380 207120 98400
rect 207380 98380 207620 98400
rect 207880 98380 208000 98400
rect 196000 98350 196100 98380
rect 196000 98150 196020 98350
rect 196090 98150 196100 98350
rect 196000 98120 196100 98150
rect 196400 98350 196600 98380
rect 196400 98150 196410 98350
rect 196480 98150 196520 98350
rect 196590 98150 196600 98350
rect 196400 98120 196600 98150
rect 196900 98350 197100 98380
rect 196900 98150 196910 98350
rect 196980 98150 197020 98350
rect 197090 98150 197100 98350
rect 196900 98120 197100 98150
rect 197400 98350 197600 98380
rect 197400 98150 197410 98350
rect 197480 98150 197520 98350
rect 197590 98150 197600 98350
rect 197400 98120 197600 98150
rect 197900 98350 198100 98380
rect 197900 98150 197910 98350
rect 197980 98150 198020 98350
rect 198090 98150 198100 98350
rect 197900 98120 198100 98150
rect 198400 98350 198600 98380
rect 198400 98150 198410 98350
rect 198480 98150 198520 98350
rect 198590 98150 198600 98350
rect 198400 98120 198600 98150
rect 198900 98350 199100 98380
rect 198900 98150 198910 98350
rect 198980 98150 199020 98350
rect 199090 98150 199100 98350
rect 198900 98120 199100 98150
rect 199400 98350 199600 98380
rect 199400 98150 199410 98350
rect 199480 98150 199520 98350
rect 199590 98150 199600 98350
rect 199400 98120 199600 98150
rect 199900 98350 200100 98380
rect 199900 98150 199910 98350
rect 199980 98150 200020 98350
rect 200090 98150 200100 98350
rect 199900 98120 200100 98150
rect 200400 98350 200600 98380
rect 200400 98150 200410 98350
rect 200480 98150 200520 98350
rect 200590 98150 200600 98350
rect 200400 98120 200600 98150
rect 200900 98350 201100 98380
rect 200900 98150 200910 98350
rect 200980 98150 201020 98350
rect 201090 98150 201100 98350
rect 200900 98120 201100 98150
rect 201400 98350 201600 98380
rect 201400 98150 201410 98350
rect 201480 98150 201520 98350
rect 201590 98150 201600 98350
rect 201400 98120 201600 98150
rect 201900 98350 202100 98380
rect 201900 98150 201910 98350
rect 201980 98150 202020 98350
rect 202090 98150 202100 98350
rect 201900 98120 202100 98150
rect 202400 98350 202600 98380
rect 202400 98150 202410 98350
rect 202480 98150 202520 98350
rect 202590 98150 202600 98350
rect 202400 98120 202600 98150
rect 202900 98350 203100 98380
rect 202900 98150 202910 98350
rect 202980 98150 203020 98350
rect 203090 98150 203100 98350
rect 202900 98120 203100 98150
rect 203400 98350 203600 98380
rect 203400 98150 203410 98350
rect 203480 98150 203520 98350
rect 203590 98150 203600 98350
rect 203400 98120 203600 98150
rect 203900 98350 204100 98380
rect 203900 98150 203910 98350
rect 203980 98150 204020 98350
rect 204090 98150 204100 98350
rect 203900 98120 204100 98150
rect 204400 98350 204600 98380
rect 204400 98150 204410 98350
rect 204480 98150 204520 98350
rect 204590 98150 204600 98350
rect 204400 98120 204600 98150
rect 204900 98350 205100 98380
rect 204900 98150 204910 98350
rect 204980 98150 205020 98350
rect 205090 98150 205100 98350
rect 204900 98120 205100 98150
rect 205400 98350 205600 98380
rect 205400 98150 205410 98350
rect 205480 98150 205520 98350
rect 205590 98150 205600 98350
rect 205400 98120 205600 98150
rect 205900 98350 206100 98380
rect 205900 98150 205910 98350
rect 205980 98150 206020 98350
rect 206090 98150 206100 98350
rect 205900 98120 206100 98150
rect 206400 98350 206600 98380
rect 206400 98150 206410 98350
rect 206480 98150 206520 98350
rect 206590 98150 206600 98350
rect 206400 98120 206600 98150
rect 206900 98350 207100 98380
rect 206900 98150 206910 98350
rect 206980 98150 207020 98350
rect 207090 98150 207100 98350
rect 206900 98120 207100 98150
rect 207400 98350 207600 98380
rect 207400 98150 207410 98350
rect 207480 98150 207520 98350
rect 207590 98150 207600 98350
rect 207400 98120 207600 98150
rect 207900 98350 208000 98380
rect 207900 98150 207910 98350
rect 207980 98150 208000 98350
rect 207900 98120 208000 98150
rect 196000 98100 196120 98120
rect 196380 98100 196620 98120
rect 196880 98100 197120 98120
rect 197380 98100 197620 98120
rect 197880 98100 198120 98120
rect 198380 98100 198620 98120
rect 198880 98100 199120 98120
rect 199380 98100 199620 98120
rect 199880 98100 200120 98120
rect 200380 98100 200620 98120
rect 200880 98100 201120 98120
rect 201380 98100 201620 98120
rect 201880 98100 202120 98120
rect 202380 98100 202620 98120
rect 202880 98100 203120 98120
rect 203380 98100 203620 98120
rect 203880 98100 204120 98120
rect 204380 98100 204620 98120
rect 204880 98100 205120 98120
rect 205380 98100 205620 98120
rect 205880 98100 206120 98120
rect 206380 98100 206620 98120
rect 206880 98100 207120 98120
rect 207380 98100 207620 98120
rect 207880 98100 208000 98120
rect 196000 98090 208000 98100
rect 196000 98020 196150 98090
rect 196350 98020 196650 98090
rect 196850 98020 197150 98090
rect 197350 98020 197650 98090
rect 197850 98020 198150 98090
rect 198350 98020 198650 98090
rect 198850 98020 199150 98090
rect 199350 98020 199650 98090
rect 199850 98020 200150 98090
rect 200350 98020 200650 98090
rect 200850 98020 201150 98090
rect 201350 98020 201650 98090
rect 201850 98020 202150 98090
rect 202350 98020 202650 98090
rect 202850 98020 203150 98090
rect 203350 98020 203650 98090
rect 203850 98020 204150 98090
rect 204350 98020 204650 98090
rect 204850 98020 205150 98090
rect 205350 98020 205650 98090
rect 205850 98020 206150 98090
rect 206350 98020 206650 98090
rect 206850 98020 207150 98090
rect 207350 98020 207650 98090
rect 207850 98020 208000 98090
rect 196000 97980 208000 98020
rect 196000 97910 196150 97980
rect 196350 97910 196650 97980
rect 196850 97910 197150 97980
rect 197350 97910 197650 97980
rect 197850 97910 198150 97980
rect 198350 97910 198650 97980
rect 198850 97910 199150 97980
rect 199350 97910 199650 97980
rect 199850 97910 200150 97980
rect 200350 97910 200650 97980
rect 200850 97910 201150 97980
rect 201350 97910 201650 97980
rect 201850 97910 202150 97980
rect 202350 97910 202650 97980
rect 202850 97910 203150 97980
rect 203350 97910 203650 97980
rect 203850 97910 204150 97980
rect 204350 97910 204650 97980
rect 204850 97910 205150 97980
rect 205350 97910 205650 97980
rect 205850 97910 206150 97980
rect 206350 97910 206650 97980
rect 206850 97910 207150 97980
rect 207350 97910 207650 97980
rect 207850 97910 208000 97980
rect 196000 97900 208000 97910
rect 196000 97880 196120 97900
rect 196380 97880 196620 97900
rect 196880 97880 197120 97900
rect 197380 97880 197620 97900
rect 197880 97880 198120 97900
rect 198380 97880 198620 97900
rect 198880 97880 199120 97900
rect 199380 97880 199620 97900
rect 199880 97880 200120 97900
rect 200380 97880 200620 97900
rect 200880 97880 201120 97900
rect 201380 97880 201620 97900
rect 201880 97880 202120 97900
rect 202380 97880 202620 97900
rect 202880 97880 203120 97900
rect 203380 97880 203620 97900
rect 203880 97880 204120 97900
rect 204380 97880 204620 97900
rect 204880 97880 205120 97900
rect 205380 97880 205620 97900
rect 205880 97880 206120 97900
rect 206380 97880 206620 97900
rect 206880 97880 207120 97900
rect 207380 97880 207620 97900
rect 207880 97880 208000 97900
rect 196000 97850 196100 97880
rect 196000 97650 196020 97850
rect 196090 97650 196100 97850
rect 196000 97620 196100 97650
rect 196400 97850 196600 97880
rect 196400 97650 196410 97850
rect 196480 97650 196520 97850
rect 196590 97650 196600 97850
rect 196400 97620 196600 97650
rect 196900 97850 197100 97880
rect 196900 97650 196910 97850
rect 196980 97650 197020 97850
rect 197090 97650 197100 97850
rect 196900 97620 197100 97650
rect 197400 97850 197600 97880
rect 197400 97650 197410 97850
rect 197480 97650 197520 97850
rect 197590 97650 197600 97850
rect 197400 97620 197600 97650
rect 197900 97850 198100 97880
rect 197900 97650 197910 97850
rect 197980 97650 198020 97850
rect 198090 97650 198100 97850
rect 197900 97620 198100 97650
rect 198400 97850 198600 97880
rect 198400 97650 198410 97850
rect 198480 97650 198520 97850
rect 198590 97650 198600 97850
rect 198400 97620 198600 97650
rect 198900 97850 199100 97880
rect 198900 97650 198910 97850
rect 198980 97650 199020 97850
rect 199090 97650 199100 97850
rect 198900 97620 199100 97650
rect 199400 97850 199600 97880
rect 199400 97650 199410 97850
rect 199480 97650 199520 97850
rect 199590 97650 199600 97850
rect 199400 97620 199600 97650
rect 199900 97850 200100 97880
rect 199900 97650 199910 97850
rect 199980 97650 200020 97850
rect 200090 97650 200100 97850
rect 199900 97620 200100 97650
rect 200400 97850 200600 97880
rect 200400 97650 200410 97850
rect 200480 97650 200520 97850
rect 200590 97650 200600 97850
rect 200400 97620 200600 97650
rect 200900 97850 201100 97880
rect 200900 97650 200910 97850
rect 200980 97650 201020 97850
rect 201090 97650 201100 97850
rect 200900 97620 201100 97650
rect 201400 97850 201600 97880
rect 201400 97650 201410 97850
rect 201480 97650 201520 97850
rect 201590 97650 201600 97850
rect 201400 97620 201600 97650
rect 201900 97850 202100 97880
rect 201900 97650 201910 97850
rect 201980 97650 202020 97850
rect 202090 97650 202100 97850
rect 201900 97620 202100 97650
rect 202400 97850 202600 97880
rect 202400 97650 202410 97850
rect 202480 97650 202520 97850
rect 202590 97650 202600 97850
rect 202400 97620 202600 97650
rect 202900 97850 203100 97880
rect 202900 97650 202910 97850
rect 202980 97650 203020 97850
rect 203090 97650 203100 97850
rect 202900 97620 203100 97650
rect 203400 97850 203600 97880
rect 203400 97650 203410 97850
rect 203480 97650 203520 97850
rect 203590 97650 203600 97850
rect 203400 97620 203600 97650
rect 203900 97850 204100 97880
rect 203900 97650 203910 97850
rect 203980 97650 204020 97850
rect 204090 97650 204100 97850
rect 203900 97620 204100 97650
rect 204400 97850 204600 97880
rect 204400 97650 204410 97850
rect 204480 97650 204520 97850
rect 204590 97650 204600 97850
rect 204400 97620 204600 97650
rect 204900 97850 205100 97880
rect 204900 97650 204910 97850
rect 204980 97650 205020 97850
rect 205090 97650 205100 97850
rect 204900 97620 205100 97650
rect 205400 97850 205600 97880
rect 205400 97650 205410 97850
rect 205480 97650 205520 97850
rect 205590 97650 205600 97850
rect 205400 97620 205600 97650
rect 205900 97850 206100 97880
rect 205900 97650 205910 97850
rect 205980 97650 206020 97850
rect 206090 97650 206100 97850
rect 205900 97620 206100 97650
rect 206400 97850 206600 97880
rect 206400 97650 206410 97850
rect 206480 97650 206520 97850
rect 206590 97650 206600 97850
rect 206400 97620 206600 97650
rect 206900 97850 207100 97880
rect 206900 97650 206910 97850
rect 206980 97650 207020 97850
rect 207090 97650 207100 97850
rect 206900 97620 207100 97650
rect 207400 97850 207600 97880
rect 207400 97650 207410 97850
rect 207480 97650 207520 97850
rect 207590 97650 207600 97850
rect 207400 97620 207600 97650
rect 207900 97850 208000 97880
rect 207900 97650 207910 97850
rect 207980 97650 208000 97850
rect 207900 97620 208000 97650
rect 196000 97600 196120 97620
rect 196380 97600 196620 97620
rect 196880 97600 197120 97620
rect 197380 97600 197620 97620
rect 197880 97600 198120 97620
rect 198380 97600 198620 97620
rect 198880 97600 199120 97620
rect 199380 97600 199620 97620
rect 199880 97600 200120 97620
rect 200380 97600 200620 97620
rect 200880 97600 201120 97620
rect 201380 97600 201620 97620
rect 201880 97600 202120 97620
rect 202380 97600 202620 97620
rect 202880 97600 203120 97620
rect 203380 97600 203620 97620
rect 203880 97600 204120 97620
rect 204380 97600 204620 97620
rect 204880 97600 205120 97620
rect 205380 97600 205620 97620
rect 205880 97600 206120 97620
rect 206380 97600 206620 97620
rect 206880 97600 207120 97620
rect 207380 97600 207620 97620
rect 207880 97600 208000 97620
rect 196000 97590 208000 97600
rect 196000 97520 196150 97590
rect 196350 97520 196650 97590
rect 196850 97520 197150 97590
rect 197350 97520 197650 97590
rect 197850 97520 198150 97590
rect 198350 97520 198650 97590
rect 198850 97520 199150 97590
rect 199350 97520 199650 97590
rect 199850 97520 200150 97590
rect 200350 97520 200650 97590
rect 200850 97520 201150 97590
rect 201350 97520 201650 97590
rect 201850 97520 202150 97590
rect 202350 97520 202650 97590
rect 202850 97520 203150 97590
rect 203350 97520 203650 97590
rect 203850 97520 204150 97590
rect 204350 97520 204650 97590
rect 204850 97520 205150 97590
rect 205350 97520 205650 97590
rect 205850 97520 206150 97590
rect 206350 97520 206650 97590
rect 206850 97520 207150 97590
rect 207350 97520 207650 97590
rect 207850 97520 208000 97590
rect 196000 97480 208000 97520
rect 196000 97410 196150 97480
rect 196350 97410 196650 97480
rect 196850 97410 197150 97480
rect 197350 97410 197650 97480
rect 197850 97410 198150 97480
rect 198350 97410 198650 97480
rect 198850 97410 199150 97480
rect 199350 97410 199650 97480
rect 199850 97410 200150 97480
rect 200350 97410 200650 97480
rect 200850 97410 201150 97480
rect 201350 97410 201650 97480
rect 201850 97410 202150 97480
rect 202350 97410 202650 97480
rect 202850 97410 203150 97480
rect 203350 97410 203650 97480
rect 203850 97410 204150 97480
rect 204350 97410 204650 97480
rect 204850 97410 205150 97480
rect 205350 97410 205650 97480
rect 205850 97410 206150 97480
rect 206350 97410 206650 97480
rect 206850 97410 207150 97480
rect 207350 97410 207650 97480
rect 207850 97410 208000 97480
rect 196000 97400 208000 97410
rect 196000 97380 196120 97400
rect 196380 97380 196620 97400
rect 196880 97380 197120 97400
rect 197380 97380 197620 97400
rect 197880 97380 198120 97400
rect 198380 97380 198620 97400
rect 198880 97380 199120 97400
rect 199380 97380 199620 97400
rect 199880 97380 200120 97400
rect 200380 97380 200620 97400
rect 200880 97380 201120 97400
rect 201380 97380 201620 97400
rect 201880 97380 202120 97400
rect 202380 97380 202620 97400
rect 202880 97380 203120 97400
rect 203380 97380 203620 97400
rect 203880 97380 204120 97400
rect 204380 97380 204620 97400
rect 204880 97380 205120 97400
rect 205380 97380 205620 97400
rect 205880 97380 206120 97400
rect 206380 97380 206620 97400
rect 206880 97380 207120 97400
rect 207380 97380 207620 97400
rect 207880 97380 208000 97400
rect 196000 97350 196100 97380
rect 196000 97150 196020 97350
rect 196090 97150 196100 97350
rect 196000 97120 196100 97150
rect 196400 97350 196600 97380
rect 196400 97150 196410 97350
rect 196480 97150 196520 97350
rect 196590 97150 196600 97350
rect 196400 97120 196600 97150
rect 196900 97350 197100 97380
rect 196900 97150 196910 97350
rect 196980 97150 197020 97350
rect 197090 97150 197100 97350
rect 196900 97120 197100 97150
rect 197400 97350 197600 97380
rect 197400 97150 197410 97350
rect 197480 97150 197520 97350
rect 197590 97150 197600 97350
rect 197400 97120 197600 97150
rect 197900 97350 198100 97380
rect 197900 97150 197910 97350
rect 197980 97150 198020 97350
rect 198090 97150 198100 97350
rect 197900 97120 198100 97150
rect 198400 97350 198600 97380
rect 198400 97150 198410 97350
rect 198480 97150 198520 97350
rect 198590 97150 198600 97350
rect 198400 97120 198600 97150
rect 198900 97350 199100 97380
rect 198900 97150 198910 97350
rect 198980 97150 199020 97350
rect 199090 97150 199100 97350
rect 198900 97120 199100 97150
rect 199400 97350 199600 97380
rect 199400 97150 199410 97350
rect 199480 97150 199520 97350
rect 199590 97150 199600 97350
rect 199400 97120 199600 97150
rect 199900 97350 200100 97380
rect 199900 97150 199910 97350
rect 199980 97150 200020 97350
rect 200090 97150 200100 97350
rect 199900 97120 200100 97150
rect 200400 97350 200600 97380
rect 200400 97150 200410 97350
rect 200480 97150 200520 97350
rect 200590 97150 200600 97350
rect 200400 97120 200600 97150
rect 200900 97350 201100 97380
rect 200900 97150 200910 97350
rect 200980 97150 201020 97350
rect 201090 97150 201100 97350
rect 200900 97120 201100 97150
rect 201400 97350 201600 97380
rect 201400 97150 201410 97350
rect 201480 97150 201520 97350
rect 201590 97150 201600 97350
rect 201400 97120 201600 97150
rect 201900 97350 202100 97380
rect 201900 97150 201910 97350
rect 201980 97150 202020 97350
rect 202090 97150 202100 97350
rect 201900 97120 202100 97150
rect 202400 97350 202600 97380
rect 202400 97150 202410 97350
rect 202480 97150 202520 97350
rect 202590 97150 202600 97350
rect 202400 97120 202600 97150
rect 202900 97350 203100 97380
rect 202900 97150 202910 97350
rect 202980 97150 203020 97350
rect 203090 97150 203100 97350
rect 202900 97120 203100 97150
rect 203400 97350 203600 97380
rect 203400 97150 203410 97350
rect 203480 97150 203520 97350
rect 203590 97150 203600 97350
rect 203400 97120 203600 97150
rect 203900 97350 204100 97380
rect 203900 97150 203910 97350
rect 203980 97150 204020 97350
rect 204090 97150 204100 97350
rect 203900 97120 204100 97150
rect 204400 97350 204600 97380
rect 204400 97150 204410 97350
rect 204480 97150 204520 97350
rect 204590 97150 204600 97350
rect 204400 97120 204600 97150
rect 204900 97350 205100 97380
rect 204900 97150 204910 97350
rect 204980 97150 205020 97350
rect 205090 97150 205100 97350
rect 204900 97120 205100 97150
rect 205400 97350 205600 97380
rect 205400 97150 205410 97350
rect 205480 97150 205520 97350
rect 205590 97150 205600 97350
rect 205400 97120 205600 97150
rect 205900 97350 206100 97380
rect 205900 97150 205910 97350
rect 205980 97150 206020 97350
rect 206090 97150 206100 97350
rect 205900 97120 206100 97150
rect 206400 97350 206600 97380
rect 206400 97150 206410 97350
rect 206480 97150 206520 97350
rect 206590 97150 206600 97350
rect 206400 97120 206600 97150
rect 206900 97350 207100 97380
rect 206900 97150 206910 97350
rect 206980 97150 207020 97350
rect 207090 97150 207100 97350
rect 206900 97120 207100 97150
rect 207400 97350 207600 97380
rect 207400 97150 207410 97350
rect 207480 97150 207520 97350
rect 207590 97150 207600 97350
rect 207400 97120 207600 97150
rect 207900 97350 208000 97380
rect 207900 97150 207910 97350
rect 207980 97150 208000 97350
rect 207900 97120 208000 97150
rect 196000 97100 196120 97120
rect 196380 97100 196620 97120
rect 196880 97100 197120 97120
rect 197380 97100 197620 97120
rect 197880 97100 198120 97120
rect 198380 97100 198620 97120
rect 198880 97100 199120 97120
rect 199380 97100 199620 97120
rect 199880 97100 200120 97120
rect 200380 97100 200620 97120
rect 200880 97100 201120 97120
rect 201380 97100 201620 97120
rect 201880 97100 202120 97120
rect 202380 97100 202620 97120
rect 202880 97100 203120 97120
rect 203380 97100 203620 97120
rect 203880 97100 204120 97120
rect 204380 97100 204620 97120
rect 204880 97100 205120 97120
rect 205380 97100 205620 97120
rect 205880 97100 206120 97120
rect 206380 97100 206620 97120
rect 206880 97100 207120 97120
rect 207380 97100 207620 97120
rect 207880 97100 208000 97120
rect 196000 97090 208000 97100
rect 196000 97020 196150 97090
rect 196350 97020 196650 97090
rect 196850 97020 197150 97090
rect 197350 97020 197650 97090
rect 197850 97020 198150 97090
rect 198350 97020 198650 97090
rect 198850 97020 199150 97090
rect 199350 97020 199650 97090
rect 199850 97020 200150 97090
rect 200350 97020 200650 97090
rect 200850 97020 201150 97090
rect 201350 97020 201650 97090
rect 201850 97020 202150 97090
rect 202350 97020 202650 97090
rect 202850 97020 203150 97090
rect 203350 97020 203650 97090
rect 203850 97020 204150 97090
rect 204350 97020 204650 97090
rect 204850 97020 205150 97090
rect 205350 97020 205650 97090
rect 205850 97020 206150 97090
rect 206350 97020 206650 97090
rect 206850 97020 207150 97090
rect 207350 97020 207650 97090
rect 207850 97020 208000 97090
rect 196000 96980 208000 97020
rect 196000 96910 196150 96980
rect 196350 96910 196650 96980
rect 196850 96910 197150 96980
rect 197350 96910 197650 96980
rect 197850 96910 198150 96980
rect 198350 96910 198650 96980
rect 198850 96910 199150 96980
rect 199350 96910 199650 96980
rect 199850 96910 200150 96980
rect 200350 96910 200650 96980
rect 200850 96910 201150 96980
rect 201350 96910 201650 96980
rect 201850 96910 202150 96980
rect 202350 96910 202650 96980
rect 202850 96910 203150 96980
rect 203350 96910 203650 96980
rect 203850 96910 204150 96980
rect 204350 96910 204650 96980
rect 204850 96910 205150 96980
rect 205350 96910 205650 96980
rect 205850 96910 206150 96980
rect 206350 96910 206650 96980
rect 206850 96910 207150 96980
rect 207350 96910 207650 96980
rect 207850 96910 208000 96980
rect 196000 96900 208000 96910
rect 196000 96880 196120 96900
rect 196380 96880 196620 96900
rect 196880 96880 197120 96900
rect 197380 96880 197620 96900
rect 197880 96880 198120 96900
rect 198380 96880 198620 96900
rect 198880 96880 199120 96900
rect 199380 96880 199620 96900
rect 199880 96880 200120 96900
rect 200380 96880 200620 96900
rect 200880 96880 201120 96900
rect 201380 96880 201620 96900
rect 201880 96880 202120 96900
rect 202380 96880 202620 96900
rect 202880 96880 203120 96900
rect 203380 96880 203620 96900
rect 203880 96880 204120 96900
rect 204380 96880 204620 96900
rect 204880 96880 205120 96900
rect 205380 96880 205620 96900
rect 205880 96880 206120 96900
rect 206380 96880 206620 96900
rect 206880 96880 207120 96900
rect 207380 96880 207620 96900
rect 207880 96880 208000 96900
rect 196000 96850 196100 96880
rect 196000 96650 196020 96850
rect 196090 96650 196100 96850
rect 196000 96620 196100 96650
rect 196400 96850 196600 96880
rect 196400 96650 196410 96850
rect 196480 96650 196520 96850
rect 196590 96650 196600 96850
rect 196400 96620 196600 96650
rect 196900 96850 197100 96880
rect 196900 96650 196910 96850
rect 196980 96650 197020 96850
rect 197090 96650 197100 96850
rect 196900 96620 197100 96650
rect 197400 96850 197600 96880
rect 197400 96650 197410 96850
rect 197480 96650 197520 96850
rect 197590 96650 197600 96850
rect 197400 96620 197600 96650
rect 197900 96850 198100 96880
rect 197900 96650 197910 96850
rect 197980 96650 198020 96850
rect 198090 96650 198100 96850
rect 197900 96620 198100 96650
rect 198400 96850 198600 96880
rect 198400 96650 198410 96850
rect 198480 96650 198520 96850
rect 198590 96650 198600 96850
rect 198400 96620 198600 96650
rect 198900 96850 199100 96880
rect 198900 96650 198910 96850
rect 198980 96650 199020 96850
rect 199090 96650 199100 96850
rect 198900 96620 199100 96650
rect 199400 96850 199600 96880
rect 199400 96650 199410 96850
rect 199480 96650 199520 96850
rect 199590 96650 199600 96850
rect 199400 96620 199600 96650
rect 199900 96850 200100 96880
rect 199900 96650 199910 96850
rect 199980 96650 200020 96850
rect 200090 96650 200100 96850
rect 199900 96620 200100 96650
rect 200400 96850 200600 96880
rect 200400 96650 200410 96850
rect 200480 96650 200520 96850
rect 200590 96650 200600 96850
rect 200400 96620 200600 96650
rect 200900 96850 201100 96880
rect 200900 96650 200910 96850
rect 200980 96650 201020 96850
rect 201090 96650 201100 96850
rect 200900 96620 201100 96650
rect 201400 96850 201600 96880
rect 201400 96650 201410 96850
rect 201480 96650 201520 96850
rect 201590 96650 201600 96850
rect 201400 96620 201600 96650
rect 201900 96850 202100 96880
rect 201900 96650 201910 96850
rect 201980 96650 202020 96850
rect 202090 96650 202100 96850
rect 201900 96620 202100 96650
rect 202400 96850 202600 96880
rect 202400 96650 202410 96850
rect 202480 96650 202520 96850
rect 202590 96650 202600 96850
rect 202400 96620 202600 96650
rect 202900 96850 203100 96880
rect 202900 96650 202910 96850
rect 202980 96650 203020 96850
rect 203090 96650 203100 96850
rect 202900 96620 203100 96650
rect 203400 96850 203600 96880
rect 203400 96650 203410 96850
rect 203480 96650 203520 96850
rect 203590 96650 203600 96850
rect 203400 96620 203600 96650
rect 203900 96850 204100 96880
rect 203900 96650 203910 96850
rect 203980 96650 204020 96850
rect 204090 96650 204100 96850
rect 203900 96620 204100 96650
rect 204400 96850 204600 96880
rect 204400 96650 204410 96850
rect 204480 96650 204520 96850
rect 204590 96650 204600 96850
rect 204400 96620 204600 96650
rect 204900 96850 205100 96880
rect 204900 96650 204910 96850
rect 204980 96650 205020 96850
rect 205090 96650 205100 96850
rect 204900 96620 205100 96650
rect 205400 96850 205600 96880
rect 205400 96650 205410 96850
rect 205480 96650 205520 96850
rect 205590 96650 205600 96850
rect 205400 96620 205600 96650
rect 205900 96850 206100 96880
rect 205900 96650 205910 96850
rect 205980 96650 206020 96850
rect 206090 96650 206100 96850
rect 205900 96620 206100 96650
rect 206400 96850 206600 96880
rect 206400 96650 206410 96850
rect 206480 96650 206520 96850
rect 206590 96650 206600 96850
rect 206400 96620 206600 96650
rect 206900 96850 207100 96880
rect 206900 96650 206910 96850
rect 206980 96650 207020 96850
rect 207090 96650 207100 96850
rect 206900 96620 207100 96650
rect 207400 96850 207600 96880
rect 207400 96650 207410 96850
rect 207480 96650 207520 96850
rect 207590 96650 207600 96850
rect 207400 96620 207600 96650
rect 207900 96850 208000 96880
rect 207900 96650 207910 96850
rect 207980 96650 208000 96850
rect 207900 96620 208000 96650
rect 196000 96600 196120 96620
rect 196380 96600 196620 96620
rect 196880 96600 197120 96620
rect 197380 96600 197620 96620
rect 197880 96600 198120 96620
rect 198380 96600 198620 96620
rect 198880 96600 199120 96620
rect 199380 96600 199620 96620
rect 199880 96600 200120 96620
rect 200380 96600 200620 96620
rect 200880 96600 201120 96620
rect 201380 96600 201620 96620
rect 201880 96600 202120 96620
rect 202380 96600 202620 96620
rect 202880 96600 203120 96620
rect 203380 96600 203620 96620
rect 203880 96600 204120 96620
rect 204380 96600 204620 96620
rect 204880 96600 205120 96620
rect 205380 96600 205620 96620
rect 205880 96600 206120 96620
rect 206380 96600 206620 96620
rect 206880 96600 207120 96620
rect 207380 96600 207620 96620
rect 207880 96600 208000 96620
rect 196000 96590 208000 96600
rect 196000 96520 196150 96590
rect 196350 96520 196650 96590
rect 196850 96520 197150 96590
rect 197350 96520 197650 96590
rect 197850 96520 198150 96590
rect 198350 96520 198650 96590
rect 198850 96520 199150 96590
rect 199350 96520 199650 96590
rect 199850 96520 200150 96590
rect 200350 96520 200650 96590
rect 200850 96520 201150 96590
rect 201350 96520 201650 96590
rect 201850 96520 202150 96590
rect 202350 96520 202650 96590
rect 202850 96520 203150 96590
rect 203350 96520 203650 96590
rect 203850 96520 204150 96590
rect 204350 96520 204650 96590
rect 204850 96520 205150 96590
rect 205350 96520 205650 96590
rect 205850 96520 206150 96590
rect 206350 96520 206650 96590
rect 206850 96520 207150 96590
rect 207350 96520 207650 96590
rect 207850 96520 208000 96590
rect 196000 96480 208000 96520
rect 196000 96410 196150 96480
rect 196350 96410 196650 96480
rect 196850 96410 197150 96480
rect 197350 96410 197650 96480
rect 197850 96410 198150 96480
rect 198350 96410 198650 96480
rect 198850 96410 199150 96480
rect 199350 96410 199650 96480
rect 199850 96410 200150 96480
rect 200350 96410 200650 96480
rect 200850 96410 201150 96480
rect 201350 96410 201650 96480
rect 201850 96410 202150 96480
rect 202350 96410 202650 96480
rect 202850 96410 203150 96480
rect 203350 96410 203650 96480
rect 203850 96410 204150 96480
rect 204350 96410 204650 96480
rect 204850 96410 205150 96480
rect 205350 96410 205650 96480
rect 205850 96410 206150 96480
rect 206350 96410 206650 96480
rect 206850 96410 207150 96480
rect 207350 96410 207650 96480
rect 207850 96410 208000 96480
rect 196000 96400 208000 96410
rect 196000 96380 196120 96400
rect 196380 96380 196620 96400
rect 196880 96380 197120 96400
rect 197380 96380 197620 96400
rect 197880 96380 198120 96400
rect 198380 96380 198620 96400
rect 198880 96380 199120 96400
rect 199380 96380 199620 96400
rect 199880 96380 200120 96400
rect 200380 96380 200620 96400
rect 200880 96380 201120 96400
rect 201380 96380 201620 96400
rect 201880 96380 202120 96400
rect 202380 96380 202620 96400
rect 202880 96380 203120 96400
rect 203380 96380 203620 96400
rect 203880 96380 204120 96400
rect 204380 96380 204620 96400
rect 204880 96380 205120 96400
rect 205380 96380 205620 96400
rect 205880 96380 206120 96400
rect 206380 96380 206620 96400
rect 206880 96380 207120 96400
rect 207380 96380 207620 96400
rect 207880 96380 208000 96400
rect 196000 96350 196100 96380
rect 196000 96150 196020 96350
rect 196090 96150 196100 96350
rect 196000 96120 196100 96150
rect 196400 96350 196600 96380
rect 196400 96150 196410 96350
rect 196480 96150 196520 96350
rect 196590 96150 196600 96350
rect 196400 96120 196600 96150
rect 196900 96350 197100 96380
rect 196900 96150 196910 96350
rect 196980 96150 197020 96350
rect 197090 96150 197100 96350
rect 196900 96120 197100 96150
rect 197400 96350 197600 96380
rect 197400 96150 197410 96350
rect 197480 96150 197520 96350
rect 197590 96150 197600 96350
rect 197400 96120 197600 96150
rect 197900 96350 198100 96380
rect 197900 96150 197910 96350
rect 197980 96150 198020 96350
rect 198090 96150 198100 96350
rect 197900 96120 198100 96150
rect 198400 96350 198600 96380
rect 198400 96150 198410 96350
rect 198480 96150 198520 96350
rect 198590 96150 198600 96350
rect 198400 96120 198600 96150
rect 198900 96350 199100 96380
rect 198900 96150 198910 96350
rect 198980 96150 199020 96350
rect 199090 96150 199100 96350
rect 198900 96120 199100 96150
rect 199400 96350 199600 96380
rect 199400 96150 199410 96350
rect 199480 96150 199520 96350
rect 199590 96150 199600 96350
rect 199400 96120 199600 96150
rect 199900 96350 200100 96380
rect 199900 96150 199910 96350
rect 199980 96150 200020 96350
rect 200090 96150 200100 96350
rect 199900 96120 200100 96150
rect 200400 96350 200600 96380
rect 200400 96150 200410 96350
rect 200480 96150 200520 96350
rect 200590 96150 200600 96350
rect 200400 96120 200600 96150
rect 200900 96350 201100 96380
rect 200900 96150 200910 96350
rect 200980 96150 201020 96350
rect 201090 96150 201100 96350
rect 200900 96120 201100 96150
rect 201400 96350 201600 96380
rect 201400 96150 201410 96350
rect 201480 96150 201520 96350
rect 201590 96150 201600 96350
rect 201400 96120 201600 96150
rect 201900 96350 202100 96380
rect 201900 96150 201910 96350
rect 201980 96150 202020 96350
rect 202090 96150 202100 96350
rect 201900 96120 202100 96150
rect 202400 96350 202600 96380
rect 202400 96150 202410 96350
rect 202480 96150 202520 96350
rect 202590 96150 202600 96350
rect 202400 96120 202600 96150
rect 202900 96350 203100 96380
rect 202900 96150 202910 96350
rect 202980 96150 203020 96350
rect 203090 96150 203100 96350
rect 202900 96120 203100 96150
rect 203400 96350 203600 96380
rect 203400 96150 203410 96350
rect 203480 96150 203520 96350
rect 203590 96150 203600 96350
rect 203400 96120 203600 96150
rect 203900 96350 204100 96380
rect 203900 96150 203910 96350
rect 203980 96150 204020 96350
rect 204090 96150 204100 96350
rect 203900 96120 204100 96150
rect 204400 96350 204600 96380
rect 204400 96150 204410 96350
rect 204480 96150 204520 96350
rect 204590 96150 204600 96350
rect 204400 96120 204600 96150
rect 204900 96350 205100 96380
rect 204900 96150 204910 96350
rect 204980 96150 205020 96350
rect 205090 96150 205100 96350
rect 204900 96120 205100 96150
rect 205400 96350 205600 96380
rect 205400 96150 205410 96350
rect 205480 96150 205520 96350
rect 205590 96150 205600 96350
rect 205400 96120 205600 96150
rect 205900 96350 206100 96380
rect 205900 96150 205910 96350
rect 205980 96150 206020 96350
rect 206090 96150 206100 96350
rect 205900 96120 206100 96150
rect 206400 96350 206600 96380
rect 206400 96150 206410 96350
rect 206480 96150 206520 96350
rect 206590 96150 206600 96350
rect 206400 96120 206600 96150
rect 206900 96350 207100 96380
rect 206900 96150 206910 96350
rect 206980 96150 207020 96350
rect 207090 96150 207100 96350
rect 206900 96120 207100 96150
rect 207400 96350 207600 96380
rect 207400 96150 207410 96350
rect 207480 96150 207520 96350
rect 207590 96150 207600 96350
rect 207400 96120 207600 96150
rect 207900 96350 208000 96380
rect 207900 96150 207910 96350
rect 207980 96150 208000 96350
rect 207900 96120 208000 96150
rect 196000 96100 196120 96120
rect 196380 96100 196620 96120
rect 196880 96100 197120 96120
rect 197380 96100 197620 96120
rect 197880 96100 198120 96120
rect 198380 96100 198620 96120
rect 198880 96100 199120 96120
rect 199380 96100 199620 96120
rect 199880 96100 200120 96120
rect 200380 96100 200620 96120
rect 200880 96100 201120 96120
rect 201380 96100 201620 96120
rect 201880 96100 202120 96120
rect 202380 96100 202620 96120
rect 202880 96100 203120 96120
rect 203380 96100 203620 96120
rect 203880 96100 204120 96120
rect 204380 96100 204620 96120
rect 204880 96100 205120 96120
rect 205380 96100 205620 96120
rect 205880 96100 206120 96120
rect 206380 96100 206620 96120
rect 206880 96100 207120 96120
rect 207380 96100 207620 96120
rect 207880 96100 208000 96120
rect 196000 96090 208000 96100
rect 196000 96020 196150 96090
rect 196350 96020 196650 96090
rect 196850 96020 197150 96090
rect 197350 96020 197650 96090
rect 197850 96020 198150 96090
rect 198350 96020 198650 96090
rect 198850 96020 199150 96090
rect 199350 96020 199650 96090
rect 199850 96020 200150 96090
rect 200350 96020 200650 96090
rect 200850 96020 201150 96090
rect 201350 96020 201650 96090
rect 201850 96020 202150 96090
rect 202350 96020 202650 96090
rect 202850 96020 203150 96090
rect 203350 96020 203650 96090
rect 203850 96020 204150 96090
rect 204350 96020 204650 96090
rect 204850 96020 205150 96090
rect 205350 96020 205650 96090
rect 205850 96020 206150 96090
rect 206350 96020 206650 96090
rect 206850 96020 207150 96090
rect 207350 96020 207650 96090
rect 207850 96020 208000 96090
rect 196000 95980 208000 96020
rect 196000 95910 196150 95980
rect 196350 95910 196650 95980
rect 196850 95910 197150 95980
rect 197350 95910 197650 95980
rect 197850 95910 198150 95980
rect 198350 95910 198650 95980
rect 198850 95910 199150 95980
rect 199350 95910 199650 95980
rect 199850 95910 200150 95980
rect 200350 95910 200650 95980
rect 200850 95910 201150 95980
rect 201350 95910 201650 95980
rect 201850 95910 202150 95980
rect 202350 95910 202650 95980
rect 202850 95910 203150 95980
rect 203350 95910 203650 95980
rect 203850 95910 204150 95980
rect 204350 95910 204650 95980
rect 204850 95910 205150 95980
rect 205350 95910 205650 95980
rect 205850 95910 206150 95980
rect 206350 95910 206650 95980
rect 206850 95910 207150 95980
rect 207350 95910 207650 95980
rect 207850 95910 208000 95980
rect 196000 95900 208000 95910
rect 196000 95880 196120 95900
rect 196380 95880 196620 95900
rect 196880 95880 197120 95900
rect 197380 95880 197620 95900
rect 197880 95880 198120 95900
rect 198380 95880 198620 95900
rect 198880 95880 199120 95900
rect 199380 95880 199620 95900
rect 199880 95880 200120 95900
rect 200380 95880 200620 95900
rect 200880 95880 201120 95900
rect 201380 95880 201620 95900
rect 201880 95880 202120 95900
rect 202380 95880 202620 95900
rect 202880 95880 203120 95900
rect 203380 95880 203620 95900
rect 203880 95880 204120 95900
rect 204380 95880 204620 95900
rect 204880 95880 205120 95900
rect 205380 95880 205620 95900
rect 205880 95880 206120 95900
rect 206380 95880 206620 95900
rect 206880 95880 207120 95900
rect 207380 95880 207620 95900
rect 207880 95880 208000 95900
rect 196000 95850 196100 95880
rect 196000 95650 196020 95850
rect 196090 95650 196100 95850
rect 196000 95620 196100 95650
rect 196400 95850 196600 95880
rect 196400 95650 196410 95850
rect 196480 95650 196520 95850
rect 196590 95650 196600 95850
rect 196400 95620 196600 95650
rect 196900 95850 197100 95880
rect 196900 95650 196910 95850
rect 196980 95650 197020 95850
rect 197090 95650 197100 95850
rect 196900 95620 197100 95650
rect 197400 95850 197600 95880
rect 197400 95650 197410 95850
rect 197480 95650 197520 95850
rect 197590 95650 197600 95850
rect 197400 95620 197600 95650
rect 197900 95850 198100 95880
rect 197900 95650 197910 95850
rect 197980 95650 198020 95850
rect 198090 95650 198100 95850
rect 197900 95620 198100 95650
rect 198400 95850 198600 95880
rect 198400 95650 198410 95850
rect 198480 95650 198520 95850
rect 198590 95650 198600 95850
rect 198400 95620 198600 95650
rect 198900 95850 199100 95880
rect 198900 95650 198910 95850
rect 198980 95650 199020 95850
rect 199090 95650 199100 95850
rect 198900 95620 199100 95650
rect 199400 95850 199600 95880
rect 199400 95650 199410 95850
rect 199480 95650 199520 95850
rect 199590 95650 199600 95850
rect 199400 95620 199600 95650
rect 199900 95850 200100 95880
rect 199900 95650 199910 95850
rect 199980 95650 200020 95850
rect 200090 95650 200100 95850
rect 199900 95620 200100 95650
rect 200400 95850 200600 95880
rect 200400 95650 200410 95850
rect 200480 95650 200520 95850
rect 200590 95650 200600 95850
rect 200400 95620 200600 95650
rect 200900 95850 201100 95880
rect 200900 95650 200910 95850
rect 200980 95650 201020 95850
rect 201090 95650 201100 95850
rect 200900 95620 201100 95650
rect 201400 95850 201600 95880
rect 201400 95650 201410 95850
rect 201480 95650 201520 95850
rect 201590 95650 201600 95850
rect 201400 95620 201600 95650
rect 201900 95850 202100 95880
rect 201900 95650 201910 95850
rect 201980 95650 202020 95850
rect 202090 95650 202100 95850
rect 201900 95620 202100 95650
rect 202400 95850 202600 95880
rect 202400 95650 202410 95850
rect 202480 95650 202520 95850
rect 202590 95650 202600 95850
rect 202400 95620 202600 95650
rect 202900 95850 203100 95880
rect 202900 95650 202910 95850
rect 202980 95650 203020 95850
rect 203090 95650 203100 95850
rect 202900 95620 203100 95650
rect 203400 95850 203600 95880
rect 203400 95650 203410 95850
rect 203480 95650 203520 95850
rect 203590 95650 203600 95850
rect 203400 95620 203600 95650
rect 203900 95850 204100 95880
rect 203900 95650 203910 95850
rect 203980 95650 204020 95850
rect 204090 95650 204100 95850
rect 203900 95620 204100 95650
rect 204400 95850 204600 95880
rect 204400 95650 204410 95850
rect 204480 95650 204520 95850
rect 204590 95650 204600 95850
rect 204400 95620 204600 95650
rect 204900 95850 205100 95880
rect 204900 95650 204910 95850
rect 204980 95650 205020 95850
rect 205090 95650 205100 95850
rect 204900 95620 205100 95650
rect 205400 95850 205600 95880
rect 205400 95650 205410 95850
rect 205480 95650 205520 95850
rect 205590 95650 205600 95850
rect 205400 95620 205600 95650
rect 205900 95850 206100 95880
rect 205900 95650 205910 95850
rect 205980 95650 206020 95850
rect 206090 95650 206100 95850
rect 205900 95620 206100 95650
rect 206400 95850 206600 95880
rect 206400 95650 206410 95850
rect 206480 95650 206520 95850
rect 206590 95650 206600 95850
rect 206400 95620 206600 95650
rect 206900 95850 207100 95880
rect 206900 95650 206910 95850
rect 206980 95650 207020 95850
rect 207090 95650 207100 95850
rect 206900 95620 207100 95650
rect 207400 95850 207600 95880
rect 207400 95650 207410 95850
rect 207480 95650 207520 95850
rect 207590 95650 207600 95850
rect 207400 95620 207600 95650
rect 207900 95850 208000 95880
rect 207900 95650 207910 95850
rect 207980 95650 208000 95850
rect 207900 95620 208000 95650
rect 196000 95600 196120 95620
rect 196380 95600 196620 95620
rect 196880 95600 197120 95620
rect 197380 95600 197620 95620
rect 197880 95600 198120 95620
rect 198380 95600 198620 95620
rect 198880 95600 199120 95620
rect 199380 95600 199620 95620
rect 199880 95600 200120 95620
rect 200380 95600 200620 95620
rect 200880 95600 201120 95620
rect 201380 95600 201620 95620
rect 201880 95600 202120 95620
rect 202380 95600 202620 95620
rect 202880 95600 203120 95620
rect 203380 95600 203620 95620
rect 203880 95600 204120 95620
rect 204380 95600 204620 95620
rect 204880 95600 205120 95620
rect 205380 95600 205620 95620
rect 205880 95600 206120 95620
rect 206380 95600 206620 95620
rect 206880 95600 207120 95620
rect 207380 95600 207620 95620
rect 207880 95600 208000 95620
rect 196000 95590 208000 95600
rect 196000 95520 196150 95590
rect 196350 95520 196650 95590
rect 196850 95520 197150 95590
rect 197350 95520 197650 95590
rect 197850 95520 198150 95590
rect 198350 95520 198650 95590
rect 198850 95520 199150 95590
rect 199350 95520 199650 95590
rect 199850 95520 200150 95590
rect 200350 95520 200650 95590
rect 200850 95520 201150 95590
rect 201350 95520 201650 95590
rect 201850 95520 202150 95590
rect 202350 95520 202650 95590
rect 202850 95520 203150 95590
rect 203350 95520 203650 95590
rect 203850 95520 204150 95590
rect 204350 95520 204650 95590
rect 204850 95520 205150 95590
rect 205350 95520 205650 95590
rect 205850 95520 206150 95590
rect 206350 95520 206650 95590
rect 206850 95520 207150 95590
rect 207350 95520 207650 95590
rect 207850 95520 208000 95590
rect 196000 95480 208000 95520
rect 196000 95410 196150 95480
rect 196350 95410 196650 95480
rect 196850 95410 197150 95480
rect 197350 95410 197650 95480
rect 197850 95410 198150 95480
rect 198350 95410 198650 95480
rect 198850 95410 199150 95480
rect 199350 95410 199650 95480
rect 199850 95410 200150 95480
rect 200350 95410 200650 95480
rect 200850 95410 201150 95480
rect 201350 95410 201650 95480
rect 201850 95410 202150 95480
rect 202350 95410 202650 95480
rect 202850 95410 203150 95480
rect 203350 95410 203650 95480
rect 203850 95410 204150 95480
rect 204350 95410 204650 95480
rect 204850 95410 205150 95480
rect 205350 95410 205650 95480
rect 205850 95410 206150 95480
rect 206350 95410 206650 95480
rect 206850 95410 207150 95480
rect 207350 95410 207650 95480
rect 207850 95410 208000 95480
rect 196000 95400 208000 95410
rect 196000 95380 196120 95400
rect 196380 95380 196620 95400
rect 196880 95380 197120 95400
rect 197380 95380 197620 95400
rect 197880 95380 198120 95400
rect 198380 95380 198620 95400
rect 198880 95380 199120 95400
rect 199380 95380 199620 95400
rect 199880 95380 200120 95400
rect 200380 95380 200620 95400
rect 200880 95380 201120 95400
rect 201380 95380 201620 95400
rect 201880 95380 202120 95400
rect 202380 95380 202620 95400
rect 202880 95380 203120 95400
rect 203380 95380 203620 95400
rect 203880 95380 204120 95400
rect 204380 95380 204620 95400
rect 204880 95380 205120 95400
rect 205380 95380 205620 95400
rect 205880 95380 206120 95400
rect 206380 95380 206620 95400
rect 206880 95380 207120 95400
rect 207380 95380 207620 95400
rect 207880 95380 208000 95400
rect 196000 95350 196100 95380
rect 196000 95150 196020 95350
rect 196090 95150 196100 95350
rect 196000 95120 196100 95150
rect 196400 95350 196600 95380
rect 196400 95150 196410 95350
rect 196480 95150 196520 95350
rect 196590 95150 196600 95350
rect 196400 95120 196600 95150
rect 196900 95350 197100 95380
rect 196900 95150 196910 95350
rect 196980 95150 197020 95350
rect 197090 95150 197100 95350
rect 196900 95120 197100 95150
rect 197400 95350 197600 95380
rect 197400 95150 197410 95350
rect 197480 95150 197520 95350
rect 197590 95150 197600 95350
rect 197400 95120 197600 95150
rect 197900 95350 198100 95380
rect 197900 95150 197910 95350
rect 197980 95150 198020 95350
rect 198090 95150 198100 95350
rect 197900 95120 198100 95150
rect 198400 95350 198600 95380
rect 198400 95150 198410 95350
rect 198480 95150 198520 95350
rect 198590 95150 198600 95350
rect 198400 95120 198600 95150
rect 198900 95350 199100 95380
rect 198900 95150 198910 95350
rect 198980 95150 199020 95350
rect 199090 95150 199100 95350
rect 198900 95120 199100 95150
rect 199400 95350 199600 95380
rect 199400 95150 199410 95350
rect 199480 95150 199520 95350
rect 199590 95150 199600 95350
rect 199400 95120 199600 95150
rect 199900 95350 200100 95380
rect 199900 95150 199910 95350
rect 199980 95150 200020 95350
rect 200090 95150 200100 95350
rect 199900 95120 200100 95150
rect 200400 95350 200600 95380
rect 200400 95150 200410 95350
rect 200480 95150 200520 95350
rect 200590 95150 200600 95350
rect 200400 95120 200600 95150
rect 200900 95350 201100 95380
rect 200900 95150 200910 95350
rect 200980 95150 201020 95350
rect 201090 95150 201100 95350
rect 200900 95120 201100 95150
rect 201400 95350 201600 95380
rect 201400 95150 201410 95350
rect 201480 95150 201520 95350
rect 201590 95150 201600 95350
rect 201400 95120 201600 95150
rect 201900 95350 202100 95380
rect 201900 95150 201910 95350
rect 201980 95150 202020 95350
rect 202090 95150 202100 95350
rect 201900 95120 202100 95150
rect 202400 95350 202600 95380
rect 202400 95150 202410 95350
rect 202480 95150 202520 95350
rect 202590 95150 202600 95350
rect 202400 95120 202600 95150
rect 202900 95350 203100 95380
rect 202900 95150 202910 95350
rect 202980 95150 203020 95350
rect 203090 95150 203100 95350
rect 202900 95120 203100 95150
rect 203400 95350 203600 95380
rect 203400 95150 203410 95350
rect 203480 95150 203520 95350
rect 203590 95150 203600 95350
rect 203400 95120 203600 95150
rect 203900 95350 204100 95380
rect 203900 95150 203910 95350
rect 203980 95150 204020 95350
rect 204090 95150 204100 95350
rect 203900 95120 204100 95150
rect 204400 95350 204600 95380
rect 204400 95150 204410 95350
rect 204480 95150 204520 95350
rect 204590 95150 204600 95350
rect 204400 95120 204600 95150
rect 204900 95350 205100 95380
rect 204900 95150 204910 95350
rect 204980 95150 205020 95350
rect 205090 95150 205100 95350
rect 204900 95120 205100 95150
rect 205400 95350 205600 95380
rect 205400 95150 205410 95350
rect 205480 95150 205520 95350
rect 205590 95150 205600 95350
rect 205400 95120 205600 95150
rect 205900 95350 206100 95380
rect 205900 95150 205910 95350
rect 205980 95150 206020 95350
rect 206090 95150 206100 95350
rect 205900 95120 206100 95150
rect 206400 95350 206600 95380
rect 206400 95150 206410 95350
rect 206480 95150 206520 95350
rect 206590 95150 206600 95350
rect 206400 95120 206600 95150
rect 206900 95350 207100 95380
rect 206900 95150 206910 95350
rect 206980 95150 207020 95350
rect 207090 95150 207100 95350
rect 206900 95120 207100 95150
rect 207400 95350 207600 95380
rect 207400 95150 207410 95350
rect 207480 95150 207520 95350
rect 207590 95150 207600 95350
rect 207400 95120 207600 95150
rect 207900 95350 208000 95380
rect 207900 95150 207910 95350
rect 207980 95150 208000 95350
rect 207900 95120 208000 95150
rect 196000 95100 196120 95120
rect 196380 95100 196620 95120
rect 196880 95100 197120 95120
rect 197380 95100 197620 95120
rect 197880 95100 198120 95120
rect 198380 95100 198620 95120
rect 198880 95100 199120 95120
rect 199380 95100 199620 95120
rect 199880 95100 200120 95120
rect 200380 95100 200620 95120
rect 200880 95100 201120 95120
rect 201380 95100 201620 95120
rect 201880 95100 202120 95120
rect 202380 95100 202620 95120
rect 202880 95100 203120 95120
rect 203380 95100 203620 95120
rect 203880 95100 204120 95120
rect 204380 95100 204620 95120
rect 204880 95100 205120 95120
rect 205380 95100 205620 95120
rect 205880 95100 206120 95120
rect 206380 95100 206620 95120
rect 206880 95100 207120 95120
rect 207380 95100 207620 95120
rect 207880 95100 208000 95120
rect 196000 95090 208000 95100
rect 196000 95020 196150 95090
rect 196350 95020 196650 95090
rect 196850 95020 197150 95090
rect 197350 95020 197650 95090
rect 197850 95020 198150 95090
rect 198350 95020 198650 95090
rect 198850 95020 199150 95090
rect 199350 95020 199650 95090
rect 199850 95020 200150 95090
rect 200350 95020 200650 95090
rect 200850 95020 201150 95090
rect 201350 95020 201650 95090
rect 201850 95020 202150 95090
rect 202350 95020 202650 95090
rect 202850 95020 203150 95090
rect 203350 95020 203650 95090
rect 203850 95020 204150 95090
rect 204350 95020 204650 95090
rect 204850 95020 205150 95090
rect 205350 95020 205650 95090
rect 205850 95020 206150 95090
rect 206350 95020 206650 95090
rect 206850 95020 207150 95090
rect 207350 95020 207650 95090
rect 207850 95020 208000 95090
rect 196000 94980 208000 95020
rect 196000 94910 196150 94980
rect 196350 94910 196650 94980
rect 196850 94910 197150 94980
rect 197350 94910 197650 94980
rect 197850 94910 198150 94980
rect 198350 94910 198650 94980
rect 198850 94910 199150 94980
rect 199350 94910 199650 94980
rect 199850 94910 200150 94980
rect 200350 94910 200650 94980
rect 200850 94910 201150 94980
rect 201350 94910 201650 94980
rect 201850 94910 202150 94980
rect 202350 94910 202650 94980
rect 202850 94910 203150 94980
rect 203350 94910 203650 94980
rect 203850 94910 204150 94980
rect 204350 94910 204650 94980
rect 204850 94910 205150 94980
rect 205350 94910 205650 94980
rect 205850 94910 206150 94980
rect 206350 94910 206650 94980
rect 206850 94910 207150 94980
rect 207350 94910 207650 94980
rect 207850 94910 208000 94980
rect 196000 94900 208000 94910
rect 196000 94880 196120 94900
rect 196380 94880 196620 94900
rect 196880 94880 197120 94900
rect 197380 94880 197620 94900
rect 197880 94880 198120 94900
rect 198380 94880 198620 94900
rect 198880 94880 199120 94900
rect 199380 94880 199620 94900
rect 199880 94880 200120 94900
rect 200380 94880 200620 94900
rect 200880 94880 201120 94900
rect 201380 94880 201620 94900
rect 201880 94880 202120 94900
rect 202380 94880 202620 94900
rect 202880 94880 203120 94900
rect 203380 94880 203620 94900
rect 203880 94880 204120 94900
rect 204380 94880 204620 94900
rect 204880 94880 205120 94900
rect 205380 94880 205620 94900
rect 205880 94880 206120 94900
rect 206380 94880 206620 94900
rect 206880 94880 207120 94900
rect 207380 94880 207620 94900
rect 207880 94880 208000 94900
rect 196000 94850 196100 94880
rect 196000 94650 196020 94850
rect 196090 94650 196100 94850
rect 196000 94620 196100 94650
rect 196400 94850 196600 94880
rect 196400 94650 196410 94850
rect 196480 94650 196520 94850
rect 196590 94650 196600 94850
rect 196400 94620 196600 94650
rect 196900 94850 197100 94880
rect 196900 94650 196910 94850
rect 196980 94650 197020 94850
rect 197090 94650 197100 94850
rect 196900 94620 197100 94650
rect 197400 94850 197600 94880
rect 197400 94650 197410 94850
rect 197480 94650 197520 94850
rect 197590 94650 197600 94850
rect 197400 94620 197600 94650
rect 197900 94850 198100 94880
rect 197900 94650 197910 94850
rect 197980 94650 198020 94850
rect 198090 94650 198100 94850
rect 197900 94620 198100 94650
rect 198400 94850 198600 94880
rect 198400 94650 198410 94850
rect 198480 94650 198520 94850
rect 198590 94650 198600 94850
rect 198400 94620 198600 94650
rect 198900 94850 199100 94880
rect 198900 94650 198910 94850
rect 198980 94650 199020 94850
rect 199090 94650 199100 94850
rect 198900 94620 199100 94650
rect 199400 94850 199600 94880
rect 199400 94650 199410 94850
rect 199480 94650 199520 94850
rect 199590 94650 199600 94850
rect 199400 94620 199600 94650
rect 199900 94850 200100 94880
rect 199900 94650 199910 94850
rect 199980 94650 200020 94850
rect 200090 94650 200100 94850
rect 199900 94620 200100 94650
rect 200400 94850 200600 94880
rect 200400 94650 200410 94850
rect 200480 94650 200520 94850
rect 200590 94650 200600 94850
rect 200400 94620 200600 94650
rect 200900 94850 201100 94880
rect 200900 94650 200910 94850
rect 200980 94650 201020 94850
rect 201090 94650 201100 94850
rect 200900 94620 201100 94650
rect 201400 94850 201600 94880
rect 201400 94650 201410 94850
rect 201480 94650 201520 94850
rect 201590 94650 201600 94850
rect 201400 94620 201600 94650
rect 201900 94850 202100 94880
rect 201900 94650 201910 94850
rect 201980 94650 202020 94850
rect 202090 94650 202100 94850
rect 201900 94620 202100 94650
rect 202400 94850 202600 94880
rect 202400 94650 202410 94850
rect 202480 94650 202520 94850
rect 202590 94650 202600 94850
rect 202400 94620 202600 94650
rect 202900 94850 203100 94880
rect 202900 94650 202910 94850
rect 202980 94650 203020 94850
rect 203090 94650 203100 94850
rect 202900 94620 203100 94650
rect 203400 94850 203600 94880
rect 203400 94650 203410 94850
rect 203480 94650 203520 94850
rect 203590 94650 203600 94850
rect 203400 94620 203600 94650
rect 203900 94850 204100 94880
rect 203900 94650 203910 94850
rect 203980 94650 204020 94850
rect 204090 94650 204100 94850
rect 203900 94620 204100 94650
rect 204400 94850 204600 94880
rect 204400 94650 204410 94850
rect 204480 94650 204520 94850
rect 204590 94650 204600 94850
rect 204400 94620 204600 94650
rect 204900 94850 205100 94880
rect 204900 94650 204910 94850
rect 204980 94650 205020 94850
rect 205090 94650 205100 94850
rect 204900 94620 205100 94650
rect 205400 94850 205600 94880
rect 205400 94650 205410 94850
rect 205480 94650 205520 94850
rect 205590 94650 205600 94850
rect 205400 94620 205600 94650
rect 205900 94850 206100 94880
rect 205900 94650 205910 94850
rect 205980 94650 206020 94850
rect 206090 94650 206100 94850
rect 205900 94620 206100 94650
rect 206400 94850 206600 94880
rect 206400 94650 206410 94850
rect 206480 94650 206520 94850
rect 206590 94650 206600 94850
rect 206400 94620 206600 94650
rect 206900 94850 207100 94880
rect 206900 94650 206910 94850
rect 206980 94650 207020 94850
rect 207090 94650 207100 94850
rect 206900 94620 207100 94650
rect 207400 94850 207600 94880
rect 207400 94650 207410 94850
rect 207480 94650 207520 94850
rect 207590 94650 207600 94850
rect 207400 94620 207600 94650
rect 207900 94850 208000 94880
rect 207900 94650 207910 94850
rect 207980 94650 208000 94850
rect 207900 94620 208000 94650
rect 196000 94600 196120 94620
rect 196380 94600 196620 94620
rect 196880 94600 197120 94620
rect 197380 94600 197620 94620
rect 197880 94600 198120 94620
rect 198380 94600 198620 94620
rect 198880 94600 199120 94620
rect 199380 94600 199620 94620
rect 199880 94600 200120 94620
rect 200380 94600 200620 94620
rect 200880 94600 201120 94620
rect 201380 94600 201620 94620
rect 201880 94600 202120 94620
rect 202380 94600 202620 94620
rect 202880 94600 203120 94620
rect 203380 94600 203620 94620
rect 203880 94600 204120 94620
rect 204380 94600 204620 94620
rect 204880 94600 205120 94620
rect 205380 94600 205620 94620
rect 205880 94600 206120 94620
rect 206380 94600 206620 94620
rect 206880 94600 207120 94620
rect 207380 94600 207620 94620
rect 207880 94600 208000 94620
rect 196000 94590 208000 94600
rect 196000 94520 196150 94590
rect 196350 94520 196650 94590
rect 196850 94520 197150 94590
rect 197350 94520 197650 94590
rect 197850 94520 198150 94590
rect 198350 94520 198650 94590
rect 198850 94520 199150 94590
rect 199350 94520 199650 94590
rect 199850 94520 200150 94590
rect 200350 94520 200650 94590
rect 200850 94520 201150 94590
rect 201350 94520 201650 94590
rect 201850 94520 202150 94590
rect 202350 94520 202650 94590
rect 202850 94520 203150 94590
rect 203350 94520 203650 94590
rect 203850 94520 204150 94590
rect 204350 94520 204650 94590
rect 204850 94520 205150 94590
rect 205350 94520 205650 94590
rect 205850 94520 206150 94590
rect 206350 94520 206650 94590
rect 206850 94520 207150 94590
rect 207350 94520 207650 94590
rect 207850 94520 208000 94590
rect 196000 94480 208000 94520
rect 196000 94410 196150 94480
rect 196350 94410 196650 94480
rect 196850 94410 197150 94480
rect 197350 94410 197650 94480
rect 197850 94410 198150 94480
rect 198350 94410 198650 94480
rect 198850 94410 199150 94480
rect 199350 94410 199650 94480
rect 199850 94410 200150 94480
rect 200350 94410 200650 94480
rect 200850 94410 201150 94480
rect 201350 94410 201650 94480
rect 201850 94410 202150 94480
rect 202350 94410 202650 94480
rect 202850 94410 203150 94480
rect 203350 94410 203650 94480
rect 203850 94410 204150 94480
rect 204350 94410 204650 94480
rect 204850 94410 205150 94480
rect 205350 94410 205650 94480
rect 205850 94410 206150 94480
rect 206350 94410 206650 94480
rect 206850 94410 207150 94480
rect 207350 94410 207650 94480
rect 207850 94410 208000 94480
rect 196000 94400 208000 94410
rect 196000 94380 196120 94400
rect 196380 94380 196620 94400
rect 196880 94380 197120 94400
rect 197380 94380 197620 94400
rect 197880 94380 198120 94400
rect 198380 94380 198620 94400
rect 198880 94380 199120 94400
rect 199380 94380 199620 94400
rect 199880 94380 200120 94400
rect 200380 94380 200620 94400
rect 200880 94380 201120 94400
rect 201380 94380 201620 94400
rect 201880 94380 202120 94400
rect 202380 94380 202620 94400
rect 202880 94380 203120 94400
rect 203380 94380 203620 94400
rect 203880 94380 204120 94400
rect 204380 94380 204620 94400
rect 204880 94380 205120 94400
rect 205380 94380 205620 94400
rect 205880 94380 206120 94400
rect 206380 94380 206620 94400
rect 206880 94380 207120 94400
rect 207380 94380 207620 94400
rect 207880 94380 208000 94400
rect 196000 94350 196100 94380
rect 196000 94150 196020 94350
rect 196090 94150 196100 94350
rect 196000 94120 196100 94150
rect 196400 94350 196600 94380
rect 196400 94150 196410 94350
rect 196480 94150 196520 94350
rect 196590 94150 196600 94350
rect 196400 94120 196600 94150
rect 196900 94350 197100 94380
rect 196900 94150 196910 94350
rect 196980 94150 197020 94350
rect 197090 94150 197100 94350
rect 196900 94120 197100 94150
rect 197400 94350 197600 94380
rect 197400 94150 197410 94350
rect 197480 94150 197520 94350
rect 197590 94150 197600 94350
rect 197400 94120 197600 94150
rect 197900 94350 198100 94380
rect 197900 94150 197910 94350
rect 197980 94150 198020 94350
rect 198090 94150 198100 94350
rect 197900 94120 198100 94150
rect 198400 94350 198600 94380
rect 198400 94150 198410 94350
rect 198480 94150 198520 94350
rect 198590 94150 198600 94350
rect 198400 94120 198600 94150
rect 198900 94350 199100 94380
rect 198900 94150 198910 94350
rect 198980 94150 199020 94350
rect 199090 94150 199100 94350
rect 198900 94120 199100 94150
rect 199400 94350 199600 94380
rect 199400 94150 199410 94350
rect 199480 94150 199520 94350
rect 199590 94150 199600 94350
rect 199400 94120 199600 94150
rect 199900 94350 200100 94380
rect 199900 94150 199910 94350
rect 199980 94150 200020 94350
rect 200090 94150 200100 94350
rect 199900 94120 200100 94150
rect 200400 94350 200600 94380
rect 200400 94150 200410 94350
rect 200480 94150 200520 94350
rect 200590 94150 200600 94350
rect 200400 94120 200600 94150
rect 200900 94350 201100 94380
rect 200900 94150 200910 94350
rect 200980 94150 201020 94350
rect 201090 94150 201100 94350
rect 200900 94120 201100 94150
rect 201400 94350 201600 94380
rect 201400 94150 201410 94350
rect 201480 94150 201520 94350
rect 201590 94150 201600 94350
rect 201400 94120 201600 94150
rect 201900 94350 202100 94380
rect 201900 94150 201910 94350
rect 201980 94150 202020 94350
rect 202090 94150 202100 94350
rect 201900 94120 202100 94150
rect 202400 94350 202600 94380
rect 202400 94150 202410 94350
rect 202480 94150 202520 94350
rect 202590 94150 202600 94350
rect 202400 94120 202600 94150
rect 202900 94350 203100 94380
rect 202900 94150 202910 94350
rect 202980 94150 203020 94350
rect 203090 94150 203100 94350
rect 202900 94120 203100 94150
rect 203400 94350 203600 94380
rect 203400 94150 203410 94350
rect 203480 94150 203520 94350
rect 203590 94150 203600 94350
rect 203400 94120 203600 94150
rect 203900 94350 204100 94380
rect 203900 94150 203910 94350
rect 203980 94150 204020 94350
rect 204090 94150 204100 94350
rect 203900 94120 204100 94150
rect 204400 94350 204600 94380
rect 204400 94150 204410 94350
rect 204480 94150 204520 94350
rect 204590 94150 204600 94350
rect 204400 94120 204600 94150
rect 204900 94350 205100 94380
rect 204900 94150 204910 94350
rect 204980 94150 205020 94350
rect 205090 94150 205100 94350
rect 204900 94120 205100 94150
rect 205400 94350 205600 94380
rect 205400 94150 205410 94350
rect 205480 94150 205520 94350
rect 205590 94150 205600 94350
rect 205400 94120 205600 94150
rect 205900 94350 206100 94380
rect 205900 94150 205910 94350
rect 205980 94150 206020 94350
rect 206090 94150 206100 94350
rect 205900 94120 206100 94150
rect 206400 94350 206600 94380
rect 206400 94150 206410 94350
rect 206480 94150 206520 94350
rect 206590 94150 206600 94350
rect 206400 94120 206600 94150
rect 206900 94350 207100 94380
rect 206900 94150 206910 94350
rect 206980 94150 207020 94350
rect 207090 94150 207100 94350
rect 206900 94120 207100 94150
rect 207400 94350 207600 94380
rect 207400 94150 207410 94350
rect 207480 94150 207520 94350
rect 207590 94150 207600 94350
rect 207400 94120 207600 94150
rect 207900 94350 208000 94380
rect 207900 94150 207910 94350
rect 207980 94150 208000 94350
rect 207900 94120 208000 94150
rect 196000 94100 196120 94120
rect 196380 94100 196620 94120
rect 196880 94100 197120 94120
rect 197380 94100 197620 94120
rect 197880 94100 198120 94120
rect 198380 94100 198620 94120
rect 198880 94100 199120 94120
rect 199380 94100 199620 94120
rect 199880 94100 200120 94120
rect 200380 94100 200620 94120
rect 200880 94100 201120 94120
rect 201380 94100 201620 94120
rect 201880 94100 202120 94120
rect 202380 94100 202620 94120
rect 202880 94100 203120 94120
rect 203380 94100 203620 94120
rect 203880 94100 204120 94120
rect 204380 94100 204620 94120
rect 204880 94100 205120 94120
rect 205380 94100 205620 94120
rect 205880 94100 206120 94120
rect 206380 94100 206620 94120
rect 206880 94100 207120 94120
rect 207380 94100 207620 94120
rect 207880 94100 208000 94120
rect 196000 94090 208000 94100
rect 196000 94020 196150 94090
rect 196350 94020 196650 94090
rect 196850 94020 197150 94090
rect 197350 94020 197650 94090
rect 197850 94020 198150 94090
rect 198350 94020 198650 94090
rect 198850 94020 199150 94090
rect 199350 94020 199650 94090
rect 199850 94020 200150 94090
rect 200350 94020 200650 94090
rect 200850 94020 201150 94090
rect 201350 94020 201650 94090
rect 201850 94020 202150 94090
rect 202350 94020 202650 94090
rect 202850 94020 203150 94090
rect 203350 94020 203650 94090
rect 203850 94020 204150 94090
rect 204350 94020 204650 94090
rect 204850 94020 205150 94090
rect 205350 94020 205650 94090
rect 205850 94020 206150 94090
rect 206350 94020 206650 94090
rect 206850 94020 207150 94090
rect 207350 94020 207650 94090
rect 207850 94020 208000 94090
rect 196000 93980 208000 94020
rect 196000 93910 196150 93980
rect 196350 93910 196650 93980
rect 196850 93910 197150 93980
rect 197350 93910 197650 93980
rect 197850 93910 198150 93980
rect 198350 93910 198650 93980
rect 198850 93910 199150 93980
rect 199350 93910 199650 93980
rect 199850 93910 200150 93980
rect 200350 93910 200650 93980
rect 200850 93910 201150 93980
rect 201350 93910 201650 93980
rect 201850 93910 202150 93980
rect 202350 93910 202650 93980
rect 202850 93910 203150 93980
rect 203350 93910 203650 93980
rect 203850 93910 204150 93980
rect 204350 93910 204650 93980
rect 204850 93910 205150 93980
rect 205350 93910 205650 93980
rect 205850 93910 206150 93980
rect 206350 93910 206650 93980
rect 206850 93910 207150 93980
rect 207350 93910 207650 93980
rect 207850 93910 208000 93980
rect 196000 93900 208000 93910
rect 196000 93880 196120 93900
rect 196380 93880 196620 93900
rect 196880 93880 197120 93900
rect 197380 93880 197620 93900
rect 197880 93880 198120 93900
rect 198380 93880 198620 93900
rect 198880 93880 199120 93900
rect 199380 93880 199620 93900
rect 199880 93880 200120 93900
rect 200380 93880 200620 93900
rect 200880 93880 201120 93900
rect 201380 93880 201620 93900
rect 201880 93880 202120 93900
rect 202380 93880 202620 93900
rect 202880 93880 203120 93900
rect 203380 93880 203620 93900
rect 203880 93880 204120 93900
rect 204380 93880 204620 93900
rect 204880 93880 205120 93900
rect 205380 93880 205620 93900
rect 205880 93880 206120 93900
rect 206380 93880 206620 93900
rect 206880 93880 207120 93900
rect 207380 93880 207620 93900
rect 207880 93880 208000 93900
rect 196000 93850 196100 93880
rect 196000 93650 196020 93850
rect 196090 93650 196100 93850
rect 196000 93620 196100 93650
rect 196400 93850 196600 93880
rect 196400 93650 196410 93850
rect 196480 93650 196520 93850
rect 196590 93650 196600 93850
rect 196400 93620 196600 93650
rect 196900 93850 197100 93880
rect 196900 93650 196910 93850
rect 196980 93650 197020 93850
rect 197090 93650 197100 93850
rect 196900 93620 197100 93650
rect 197400 93850 197600 93880
rect 197400 93650 197410 93850
rect 197480 93650 197520 93850
rect 197590 93650 197600 93850
rect 197400 93620 197600 93650
rect 197900 93850 198100 93880
rect 197900 93650 197910 93850
rect 197980 93650 198020 93850
rect 198090 93650 198100 93850
rect 197900 93620 198100 93650
rect 198400 93850 198600 93880
rect 198400 93650 198410 93850
rect 198480 93650 198520 93850
rect 198590 93650 198600 93850
rect 198400 93620 198600 93650
rect 198900 93850 199100 93880
rect 198900 93650 198910 93850
rect 198980 93650 199020 93850
rect 199090 93650 199100 93850
rect 198900 93620 199100 93650
rect 199400 93850 199600 93880
rect 199400 93650 199410 93850
rect 199480 93650 199520 93850
rect 199590 93650 199600 93850
rect 199400 93620 199600 93650
rect 199900 93850 200100 93880
rect 199900 93650 199910 93850
rect 199980 93650 200020 93850
rect 200090 93650 200100 93850
rect 199900 93620 200100 93650
rect 200400 93850 200600 93880
rect 200400 93650 200410 93850
rect 200480 93650 200520 93850
rect 200590 93650 200600 93850
rect 200400 93620 200600 93650
rect 200900 93850 201100 93880
rect 200900 93650 200910 93850
rect 200980 93650 201020 93850
rect 201090 93650 201100 93850
rect 200900 93620 201100 93650
rect 201400 93850 201600 93880
rect 201400 93650 201410 93850
rect 201480 93650 201520 93850
rect 201590 93650 201600 93850
rect 201400 93620 201600 93650
rect 201900 93850 202100 93880
rect 201900 93650 201910 93850
rect 201980 93650 202020 93850
rect 202090 93650 202100 93850
rect 201900 93620 202100 93650
rect 202400 93850 202600 93880
rect 202400 93650 202410 93850
rect 202480 93650 202520 93850
rect 202590 93650 202600 93850
rect 202400 93620 202600 93650
rect 202900 93850 203100 93880
rect 202900 93650 202910 93850
rect 202980 93650 203020 93850
rect 203090 93650 203100 93850
rect 202900 93620 203100 93650
rect 203400 93850 203600 93880
rect 203400 93650 203410 93850
rect 203480 93650 203520 93850
rect 203590 93650 203600 93850
rect 203400 93620 203600 93650
rect 203900 93850 204100 93880
rect 203900 93650 203910 93850
rect 203980 93650 204020 93850
rect 204090 93650 204100 93850
rect 203900 93620 204100 93650
rect 204400 93850 204600 93880
rect 204400 93650 204410 93850
rect 204480 93650 204520 93850
rect 204590 93650 204600 93850
rect 204400 93620 204600 93650
rect 204900 93850 205100 93880
rect 204900 93650 204910 93850
rect 204980 93650 205020 93850
rect 205090 93650 205100 93850
rect 204900 93620 205100 93650
rect 205400 93850 205600 93880
rect 205400 93650 205410 93850
rect 205480 93650 205520 93850
rect 205590 93650 205600 93850
rect 205400 93620 205600 93650
rect 205900 93850 206100 93880
rect 205900 93650 205910 93850
rect 205980 93650 206020 93850
rect 206090 93650 206100 93850
rect 205900 93620 206100 93650
rect 206400 93850 206600 93880
rect 206400 93650 206410 93850
rect 206480 93650 206520 93850
rect 206590 93650 206600 93850
rect 206400 93620 206600 93650
rect 206900 93850 207100 93880
rect 206900 93650 206910 93850
rect 206980 93650 207020 93850
rect 207090 93650 207100 93850
rect 206900 93620 207100 93650
rect 207400 93850 207600 93880
rect 207400 93650 207410 93850
rect 207480 93650 207520 93850
rect 207590 93650 207600 93850
rect 207400 93620 207600 93650
rect 207900 93850 208000 93880
rect 207900 93650 207910 93850
rect 207980 93650 208000 93850
rect 207900 93620 208000 93650
rect 196000 93600 196120 93620
rect 196380 93600 196620 93620
rect 196880 93600 197120 93620
rect 197380 93600 197620 93620
rect 197880 93600 198120 93620
rect 198380 93600 198620 93620
rect 198880 93600 199120 93620
rect 199380 93600 199620 93620
rect 199880 93600 200120 93620
rect 200380 93600 200620 93620
rect 200880 93600 201120 93620
rect 201380 93600 201620 93620
rect 201880 93600 202120 93620
rect 202380 93600 202620 93620
rect 202880 93600 203120 93620
rect 203380 93600 203620 93620
rect 203880 93600 204120 93620
rect 204380 93600 204620 93620
rect 204880 93600 205120 93620
rect 205380 93600 205620 93620
rect 205880 93600 206120 93620
rect 206380 93600 206620 93620
rect 206880 93600 207120 93620
rect 207380 93600 207620 93620
rect 207880 93600 208000 93620
rect 196000 93590 208000 93600
rect 196000 93520 196150 93590
rect 196350 93520 196650 93590
rect 196850 93520 197150 93590
rect 197350 93520 197650 93590
rect 197850 93520 198150 93590
rect 198350 93520 198650 93590
rect 198850 93520 199150 93590
rect 199350 93520 199650 93590
rect 199850 93520 200150 93590
rect 200350 93520 200650 93590
rect 200850 93520 201150 93590
rect 201350 93520 201650 93590
rect 201850 93520 202150 93590
rect 202350 93520 202650 93590
rect 202850 93520 203150 93590
rect 203350 93520 203650 93590
rect 203850 93520 204150 93590
rect 204350 93520 204650 93590
rect 204850 93520 205150 93590
rect 205350 93520 205650 93590
rect 205850 93520 206150 93590
rect 206350 93520 206650 93590
rect 206850 93520 207150 93590
rect 207350 93520 207650 93590
rect 207850 93520 208000 93590
rect 196000 93480 208000 93520
rect 196000 93410 196150 93480
rect 196350 93410 196650 93480
rect 196850 93410 197150 93480
rect 197350 93410 197650 93480
rect 197850 93410 198150 93480
rect 198350 93410 198650 93480
rect 198850 93410 199150 93480
rect 199350 93410 199650 93480
rect 199850 93410 200150 93480
rect 200350 93410 200650 93480
rect 200850 93410 201150 93480
rect 201350 93410 201650 93480
rect 201850 93410 202150 93480
rect 202350 93410 202650 93480
rect 202850 93410 203150 93480
rect 203350 93410 203650 93480
rect 203850 93410 204150 93480
rect 204350 93410 204650 93480
rect 204850 93410 205150 93480
rect 205350 93410 205650 93480
rect 205850 93410 206150 93480
rect 206350 93410 206650 93480
rect 206850 93410 207150 93480
rect 207350 93410 207650 93480
rect 207850 93410 208000 93480
rect 196000 93400 208000 93410
rect 196000 93380 196120 93400
rect 196380 93380 196620 93400
rect 196880 93380 197120 93400
rect 197380 93380 197620 93400
rect 197880 93380 198120 93400
rect 198380 93380 198620 93400
rect 198880 93380 199120 93400
rect 199380 93380 199620 93400
rect 199880 93380 200120 93400
rect 200380 93380 200620 93400
rect 200880 93380 201120 93400
rect 201380 93380 201620 93400
rect 201880 93380 202120 93400
rect 202380 93380 202620 93400
rect 202880 93380 203120 93400
rect 203380 93380 203620 93400
rect 203880 93380 204120 93400
rect 204380 93380 204620 93400
rect 204880 93380 205120 93400
rect 205380 93380 205620 93400
rect 205880 93380 206120 93400
rect 206380 93380 206620 93400
rect 206880 93380 207120 93400
rect 207380 93380 207620 93400
rect 207880 93380 208000 93400
rect 196000 93350 196100 93380
rect 196000 93150 196020 93350
rect 196090 93150 196100 93350
rect 196000 93120 196100 93150
rect 196400 93350 196600 93380
rect 196400 93150 196410 93350
rect 196480 93150 196520 93350
rect 196590 93150 196600 93350
rect 196400 93120 196600 93150
rect 196900 93350 197100 93380
rect 196900 93150 196910 93350
rect 196980 93150 197020 93350
rect 197090 93150 197100 93350
rect 196900 93120 197100 93150
rect 197400 93350 197600 93380
rect 197400 93150 197410 93350
rect 197480 93150 197520 93350
rect 197590 93150 197600 93350
rect 197400 93120 197600 93150
rect 197900 93350 198100 93380
rect 197900 93150 197910 93350
rect 197980 93150 198020 93350
rect 198090 93150 198100 93350
rect 197900 93120 198100 93150
rect 198400 93350 198600 93380
rect 198400 93150 198410 93350
rect 198480 93150 198520 93350
rect 198590 93150 198600 93350
rect 198400 93120 198600 93150
rect 198900 93350 199100 93380
rect 198900 93150 198910 93350
rect 198980 93150 199020 93350
rect 199090 93150 199100 93350
rect 198900 93120 199100 93150
rect 199400 93350 199600 93380
rect 199400 93150 199410 93350
rect 199480 93150 199520 93350
rect 199590 93150 199600 93350
rect 199400 93120 199600 93150
rect 199900 93350 200100 93380
rect 199900 93150 199910 93350
rect 199980 93150 200020 93350
rect 200090 93150 200100 93350
rect 199900 93120 200100 93150
rect 200400 93350 200600 93380
rect 200400 93150 200410 93350
rect 200480 93150 200520 93350
rect 200590 93150 200600 93350
rect 200400 93120 200600 93150
rect 200900 93350 201100 93380
rect 200900 93150 200910 93350
rect 200980 93150 201020 93350
rect 201090 93150 201100 93350
rect 200900 93120 201100 93150
rect 201400 93350 201600 93380
rect 201400 93150 201410 93350
rect 201480 93150 201520 93350
rect 201590 93150 201600 93350
rect 201400 93120 201600 93150
rect 201900 93350 202100 93380
rect 201900 93150 201910 93350
rect 201980 93150 202020 93350
rect 202090 93150 202100 93350
rect 201900 93120 202100 93150
rect 202400 93350 202600 93380
rect 202400 93150 202410 93350
rect 202480 93150 202520 93350
rect 202590 93150 202600 93350
rect 202400 93120 202600 93150
rect 202900 93350 203100 93380
rect 202900 93150 202910 93350
rect 202980 93150 203020 93350
rect 203090 93150 203100 93350
rect 202900 93120 203100 93150
rect 203400 93350 203600 93380
rect 203400 93150 203410 93350
rect 203480 93150 203520 93350
rect 203590 93150 203600 93350
rect 203400 93120 203600 93150
rect 203900 93350 204100 93380
rect 203900 93150 203910 93350
rect 203980 93150 204020 93350
rect 204090 93150 204100 93350
rect 203900 93120 204100 93150
rect 204400 93350 204600 93380
rect 204400 93150 204410 93350
rect 204480 93150 204520 93350
rect 204590 93150 204600 93350
rect 204400 93120 204600 93150
rect 204900 93350 205100 93380
rect 204900 93150 204910 93350
rect 204980 93150 205020 93350
rect 205090 93150 205100 93350
rect 204900 93120 205100 93150
rect 205400 93350 205600 93380
rect 205400 93150 205410 93350
rect 205480 93150 205520 93350
rect 205590 93150 205600 93350
rect 205400 93120 205600 93150
rect 205900 93350 206100 93380
rect 205900 93150 205910 93350
rect 205980 93150 206020 93350
rect 206090 93150 206100 93350
rect 205900 93120 206100 93150
rect 206400 93350 206600 93380
rect 206400 93150 206410 93350
rect 206480 93150 206520 93350
rect 206590 93150 206600 93350
rect 206400 93120 206600 93150
rect 206900 93350 207100 93380
rect 206900 93150 206910 93350
rect 206980 93150 207020 93350
rect 207090 93150 207100 93350
rect 206900 93120 207100 93150
rect 207400 93350 207600 93380
rect 207400 93150 207410 93350
rect 207480 93150 207520 93350
rect 207590 93150 207600 93350
rect 207400 93120 207600 93150
rect 207900 93350 208000 93380
rect 207900 93150 207910 93350
rect 207980 93150 208000 93350
rect 207900 93120 208000 93150
rect 196000 93100 196120 93120
rect 196380 93100 196620 93120
rect 196880 93100 197120 93120
rect 197380 93100 197620 93120
rect 197880 93100 198120 93120
rect 198380 93100 198620 93120
rect 198880 93100 199120 93120
rect 199380 93100 199620 93120
rect 199880 93100 200120 93120
rect 200380 93100 200620 93120
rect 200880 93100 201120 93120
rect 201380 93100 201620 93120
rect 201880 93100 202120 93120
rect 202380 93100 202620 93120
rect 202880 93100 203120 93120
rect 203380 93100 203620 93120
rect 203880 93100 204120 93120
rect 204380 93100 204620 93120
rect 204880 93100 205120 93120
rect 205380 93100 205620 93120
rect 205880 93100 206120 93120
rect 206380 93100 206620 93120
rect 206880 93100 207120 93120
rect 207380 93100 207620 93120
rect 207880 93100 208000 93120
rect 196000 93090 208000 93100
rect 196000 93020 196150 93090
rect 196350 93020 196650 93090
rect 196850 93020 197150 93090
rect 197350 93020 197650 93090
rect 197850 93020 198150 93090
rect 198350 93020 198650 93090
rect 198850 93020 199150 93090
rect 199350 93020 199650 93090
rect 199850 93020 200150 93090
rect 200350 93020 200650 93090
rect 200850 93020 201150 93090
rect 201350 93020 201650 93090
rect 201850 93020 202150 93090
rect 202350 93020 202650 93090
rect 202850 93020 203150 93090
rect 203350 93020 203650 93090
rect 203850 93020 204150 93090
rect 204350 93020 204650 93090
rect 204850 93020 205150 93090
rect 205350 93020 205650 93090
rect 205850 93020 206150 93090
rect 206350 93020 206650 93090
rect 206850 93020 207150 93090
rect 207350 93020 207650 93090
rect 207850 93020 208000 93090
rect 196000 92980 208000 93020
rect 196000 92910 196150 92980
rect 196350 92910 196650 92980
rect 196850 92910 197150 92980
rect 197350 92910 197650 92980
rect 197850 92910 198150 92980
rect 198350 92910 198650 92980
rect 198850 92910 199150 92980
rect 199350 92910 199650 92980
rect 199850 92910 200150 92980
rect 200350 92910 200650 92980
rect 200850 92910 201150 92980
rect 201350 92910 201650 92980
rect 201850 92910 202150 92980
rect 202350 92910 202650 92980
rect 202850 92910 203150 92980
rect 203350 92910 203650 92980
rect 203850 92910 204150 92980
rect 204350 92910 204650 92980
rect 204850 92910 205150 92980
rect 205350 92910 205650 92980
rect 205850 92910 206150 92980
rect 206350 92910 206650 92980
rect 206850 92910 207150 92980
rect 207350 92910 207650 92980
rect 207850 92910 208000 92980
rect 196000 92900 208000 92910
rect 196000 92880 196120 92900
rect 196380 92880 196620 92900
rect 196880 92880 197120 92900
rect 197380 92880 197620 92900
rect 197880 92880 198120 92900
rect 198380 92880 198620 92900
rect 198880 92880 199120 92900
rect 199380 92880 199620 92900
rect 199880 92880 200120 92900
rect 200380 92880 200620 92900
rect 200880 92880 201120 92900
rect 201380 92880 201620 92900
rect 201880 92880 202120 92900
rect 202380 92880 202620 92900
rect 202880 92880 203120 92900
rect 203380 92880 203620 92900
rect 203880 92880 204120 92900
rect 204380 92880 204620 92900
rect 204880 92880 205120 92900
rect 205380 92880 205620 92900
rect 205880 92880 206120 92900
rect 206380 92880 206620 92900
rect 206880 92880 207120 92900
rect 207380 92880 207620 92900
rect 207880 92880 208000 92900
rect 196000 92850 196100 92880
rect 196000 92650 196020 92850
rect 196090 92650 196100 92850
rect 196000 92620 196100 92650
rect 196400 92850 196600 92880
rect 196400 92650 196410 92850
rect 196480 92650 196520 92850
rect 196590 92650 196600 92850
rect 196400 92620 196600 92650
rect 196900 92850 197100 92880
rect 196900 92650 196910 92850
rect 196980 92650 197020 92850
rect 197090 92650 197100 92850
rect 196900 92620 197100 92650
rect 197400 92850 197600 92880
rect 197400 92650 197410 92850
rect 197480 92650 197520 92850
rect 197590 92650 197600 92850
rect 197400 92620 197600 92650
rect 197900 92850 198100 92880
rect 197900 92650 197910 92850
rect 197980 92650 198020 92850
rect 198090 92650 198100 92850
rect 197900 92620 198100 92650
rect 198400 92850 198600 92880
rect 198400 92650 198410 92850
rect 198480 92650 198520 92850
rect 198590 92650 198600 92850
rect 198400 92620 198600 92650
rect 198900 92850 199100 92880
rect 198900 92650 198910 92850
rect 198980 92650 199020 92850
rect 199090 92650 199100 92850
rect 198900 92620 199100 92650
rect 199400 92850 199600 92880
rect 199400 92650 199410 92850
rect 199480 92650 199520 92850
rect 199590 92650 199600 92850
rect 199400 92620 199600 92650
rect 199900 92850 200100 92880
rect 199900 92650 199910 92850
rect 199980 92650 200020 92850
rect 200090 92650 200100 92850
rect 199900 92620 200100 92650
rect 200400 92850 200600 92880
rect 200400 92650 200410 92850
rect 200480 92650 200520 92850
rect 200590 92650 200600 92850
rect 200400 92620 200600 92650
rect 200900 92850 201100 92880
rect 200900 92650 200910 92850
rect 200980 92650 201020 92850
rect 201090 92650 201100 92850
rect 200900 92620 201100 92650
rect 201400 92850 201600 92880
rect 201400 92650 201410 92850
rect 201480 92650 201520 92850
rect 201590 92650 201600 92850
rect 201400 92620 201600 92650
rect 201900 92850 202100 92880
rect 201900 92650 201910 92850
rect 201980 92650 202020 92850
rect 202090 92650 202100 92850
rect 201900 92620 202100 92650
rect 202400 92850 202600 92880
rect 202400 92650 202410 92850
rect 202480 92650 202520 92850
rect 202590 92650 202600 92850
rect 202400 92620 202600 92650
rect 202900 92850 203100 92880
rect 202900 92650 202910 92850
rect 202980 92650 203020 92850
rect 203090 92650 203100 92850
rect 202900 92620 203100 92650
rect 203400 92850 203600 92880
rect 203400 92650 203410 92850
rect 203480 92650 203520 92850
rect 203590 92650 203600 92850
rect 203400 92620 203600 92650
rect 203900 92850 204100 92880
rect 203900 92650 203910 92850
rect 203980 92650 204020 92850
rect 204090 92650 204100 92850
rect 203900 92620 204100 92650
rect 204400 92850 204600 92880
rect 204400 92650 204410 92850
rect 204480 92650 204520 92850
rect 204590 92650 204600 92850
rect 204400 92620 204600 92650
rect 204900 92850 205100 92880
rect 204900 92650 204910 92850
rect 204980 92650 205020 92850
rect 205090 92650 205100 92850
rect 204900 92620 205100 92650
rect 205400 92850 205600 92880
rect 205400 92650 205410 92850
rect 205480 92650 205520 92850
rect 205590 92650 205600 92850
rect 205400 92620 205600 92650
rect 205900 92850 206100 92880
rect 205900 92650 205910 92850
rect 205980 92650 206020 92850
rect 206090 92650 206100 92850
rect 205900 92620 206100 92650
rect 206400 92850 206600 92880
rect 206400 92650 206410 92850
rect 206480 92650 206520 92850
rect 206590 92650 206600 92850
rect 206400 92620 206600 92650
rect 206900 92850 207100 92880
rect 206900 92650 206910 92850
rect 206980 92650 207020 92850
rect 207090 92650 207100 92850
rect 206900 92620 207100 92650
rect 207400 92850 207600 92880
rect 207400 92650 207410 92850
rect 207480 92650 207520 92850
rect 207590 92650 207600 92850
rect 207400 92620 207600 92650
rect 207900 92850 208000 92880
rect 207900 92650 207910 92850
rect 207980 92650 208000 92850
rect 207900 92620 208000 92650
rect 196000 92600 196120 92620
rect 196380 92600 196620 92620
rect 196880 92600 197120 92620
rect 197380 92600 197620 92620
rect 197880 92600 198120 92620
rect 198380 92600 198620 92620
rect 198880 92600 199120 92620
rect 199380 92600 199620 92620
rect 199880 92600 200120 92620
rect 200380 92600 200620 92620
rect 200880 92600 201120 92620
rect 201380 92600 201620 92620
rect 201880 92600 202120 92620
rect 202380 92600 202620 92620
rect 202880 92600 203120 92620
rect 203380 92600 203620 92620
rect 203880 92600 204120 92620
rect 204380 92600 204620 92620
rect 204880 92600 205120 92620
rect 205380 92600 205620 92620
rect 205880 92600 206120 92620
rect 206380 92600 206620 92620
rect 206880 92600 207120 92620
rect 207380 92600 207620 92620
rect 207880 92600 208000 92620
rect 196000 92590 208000 92600
rect 196000 92520 196150 92590
rect 196350 92520 196650 92590
rect 196850 92520 197150 92590
rect 197350 92520 197650 92590
rect 197850 92520 198150 92590
rect 198350 92520 198650 92590
rect 198850 92520 199150 92590
rect 199350 92520 199650 92590
rect 199850 92520 200150 92590
rect 200350 92520 200650 92590
rect 200850 92520 201150 92590
rect 201350 92520 201650 92590
rect 201850 92520 202150 92590
rect 202350 92520 202650 92590
rect 202850 92520 203150 92590
rect 203350 92520 203650 92590
rect 203850 92520 204150 92590
rect 204350 92520 204650 92590
rect 204850 92520 205150 92590
rect 205350 92520 205650 92590
rect 205850 92520 206150 92590
rect 206350 92520 206650 92590
rect 206850 92520 207150 92590
rect 207350 92520 207650 92590
rect 207850 92520 208000 92590
rect 196000 92480 208000 92520
rect 196000 92410 196150 92480
rect 196350 92410 196650 92480
rect 196850 92410 197150 92480
rect 197350 92410 197650 92480
rect 197850 92410 198150 92480
rect 198350 92410 198650 92480
rect 198850 92410 199150 92480
rect 199350 92410 199650 92480
rect 199850 92410 200150 92480
rect 200350 92410 200650 92480
rect 200850 92410 201150 92480
rect 201350 92410 201650 92480
rect 201850 92410 202150 92480
rect 202350 92410 202650 92480
rect 202850 92410 203150 92480
rect 203350 92410 203650 92480
rect 203850 92410 204150 92480
rect 204350 92410 204650 92480
rect 204850 92410 205150 92480
rect 205350 92410 205650 92480
rect 205850 92410 206150 92480
rect 206350 92410 206650 92480
rect 206850 92410 207150 92480
rect 207350 92410 207650 92480
rect 207850 92410 208000 92480
rect 196000 92400 208000 92410
rect 196000 92380 196120 92400
rect 196380 92380 196620 92400
rect 196880 92380 197120 92400
rect 197380 92380 197620 92400
rect 197880 92380 198120 92400
rect 198380 92380 198620 92400
rect 198880 92380 199120 92400
rect 199380 92380 199620 92400
rect 199880 92380 200120 92400
rect 200380 92380 200620 92400
rect 200880 92380 201120 92400
rect 201380 92380 201620 92400
rect 201880 92380 202120 92400
rect 202380 92380 202620 92400
rect 202880 92380 203120 92400
rect 203380 92380 203620 92400
rect 203880 92380 204120 92400
rect 204380 92380 204620 92400
rect 204880 92380 205120 92400
rect 205380 92380 205620 92400
rect 205880 92380 206120 92400
rect 206380 92380 206620 92400
rect 206880 92380 207120 92400
rect 207380 92380 207620 92400
rect 207880 92380 208000 92400
rect 196000 92350 196100 92380
rect 196000 92150 196020 92350
rect 196090 92150 196100 92350
rect 196000 92120 196100 92150
rect 196400 92350 196600 92380
rect 196400 92150 196410 92350
rect 196480 92150 196520 92350
rect 196590 92150 196600 92350
rect 196400 92120 196600 92150
rect 196900 92350 197100 92380
rect 196900 92150 196910 92350
rect 196980 92150 197020 92350
rect 197090 92150 197100 92350
rect 196900 92120 197100 92150
rect 197400 92350 197600 92380
rect 197400 92150 197410 92350
rect 197480 92150 197520 92350
rect 197590 92150 197600 92350
rect 197400 92120 197600 92150
rect 197900 92350 198100 92380
rect 197900 92150 197910 92350
rect 197980 92150 198020 92350
rect 198090 92150 198100 92350
rect 197900 92120 198100 92150
rect 198400 92350 198600 92380
rect 198400 92150 198410 92350
rect 198480 92150 198520 92350
rect 198590 92150 198600 92350
rect 198400 92120 198600 92150
rect 198900 92350 199100 92380
rect 198900 92150 198910 92350
rect 198980 92150 199020 92350
rect 199090 92150 199100 92350
rect 198900 92120 199100 92150
rect 199400 92350 199600 92380
rect 199400 92150 199410 92350
rect 199480 92150 199520 92350
rect 199590 92150 199600 92350
rect 199400 92120 199600 92150
rect 199900 92350 200100 92380
rect 199900 92150 199910 92350
rect 199980 92150 200020 92350
rect 200090 92150 200100 92350
rect 199900 92120 200100 92150
rect 200400 92350 200600 92380
rect 200400 92150 200410 92350
rect 200480 92150 200520 92350
rect 200590 92150 200600 92350
rect 200400 92120 200600 92150
rect 200900 92350 201100 92380
rect 200900 92150 200910 92350
rect 200980 92150 201020 92350
rect 201090 92150 201100 92350
rect 200900 92120 201100 92150
rect 201400 92350 201600 92380
rect 201400 92150 201410 92350
rect 201480 92150 201520 92350
rect 201590 92150 201600 92350
rect 201400 92120 201600 92150
rect 201900 92350 202100 92380
rect 201900 92150 201910 92350
rect 201980 92150 202020 92350
rect 202090 92150 202100 92350
rect 201900 92120 202100 92150
rect 202400 92350 202600 92380
rect 202400 92150 202410 92350
rect 202480 92150 202520 92350
rect 202590 92150 202600 92350
rect 202400 92120 202600 92150
rect 202900 92350 203100 92380
rect 202900 92150 202910 92350
rect 202980 92150 203020 92350
rect 203090 92150 203100 92350
rect 202900 92120 203100 92150
rect 203400 92350 203600 92380
rect 203400 92150 203410 92350
rect 203480 92150 203520 92350
rect 203590 92150 203600 92350
rect 203400 92120 203600 92150
rect 203900 92350 204100 92380
rect 203900 92150 203910 92350
rect 203980 92150 204020 92350
rect 204090 92150 204100 92350
rect 203900 92120 204100 92150
rect 204400 92350 204600 92380
rect 204400 92150 204410 92350
rect 204480 92150 204520 92350
rect 204590 92150 204600 92350
rect 204400 92120 204600 92150
rect 204900 92350 205100 92380
rect 204900 92150 204910 92350
rect 204980 92150 205020 92350
rect 205090 92150 205100 92350
rect 204900 92120 205100 92150
rect 205400 92350 205600 92380
rect 205400 92150 205410 92350
rect 205480 92150 205520 92350
rect 205590 92150 205600 92350
rect 205400 92120 205600 92150
rect 205900 92350 206100 92380
rect 205900 92150 205910 92350
rect 205980 92150 206020 92350
rect 206090 92150 206100 92350
rect 205900 92120 206100 92150
rect 206400 92350 206600 92380
rect 206400 92150 206410 92350
rect 206480 92150 206520 92350
rect 206590 92150 206600 92350
rect 206400 92120 206600 92150
rect 206900 92350 207100 92380
rect 206900 92150 206910 92350
rect 206980 92150 207020 92350
rect 207090 92150 207100 92350
rect 206900 92120 207100 92150
rect 207400 92350 207600 92380
rect 207400 92150 207410 92350
rect 207480 92150 207520 92350
rect 207590 92150 207600 92350
rect 207400 92120 207600 92150
rect 207900 92350 208000 92380
rect 207900 92150 207910 92350
rect 207980 92150 208000 92350
rect 207900 92120 208000 92150
rect 196000 92100 196120 92120
rect 196380 92100 196620 92120
rect 196880 92100 197120 92120
rect 197380 92100 197620 92120
rect 197880 92100 198120 92120
rect 198380 92100 198620 92120
rect 198880 92100 199120 92120
rect 199380 92100 199620 92120
rect 199880 92100 200120 92120
rect 200380 92100 200620 92120
rect 200880 92100 201120 92120
rect 201380 92100 201620 92120
rect 201880 92100 202120 92120
rect 202380 92100 202620 92120
rect 202880 92100 203120 92120
rect 203380 92100 203620 92120
rect 203880 92100 204120 92120
rect 204380 92100 204620 92120
rect 204880 92100 205120 92120
rect 205380 92100 205620 92120
rect 205880 92100 206120 92120
rect 206380 92100 206620 92120
rect 206880 92100 207120 92120
rect 207380 92100 207620 92120
rect 207880 92100 208000 92120
rect 196000 92090 208000 92100
rect 196000 92020 196150 92090
rect 196350 92020 196650 92090
rect 196850 92020 197150 92090
rect 197350 92020 197650 92090
rect 197850 92020 198150 92090
rect 198350 92020 198650 92090
rect 198850 92020 199150 92090
rect 199350 92020 199650 92090
rect 199850 92020 200150 92090
rect 200350 92020 200650 92090
rect 200850 92020 201150 92090
rect 201350 92020 201650 92090
rect 201850 92020 202150 92090
rect 202350 92020 202650 92090
rect 202850 92020 203150 92090
rect 203350 92020 203650 92090
rect 203850 92020 204150 92090
rect 204350 92020 204650 92090
rect 204850 92020 205150 92090
rect 205350 92020 205650 92090
rect 205850 92020 206150 92090
rect 206350 92020 206650 92090
rect 206850 92020 207150 92090
rect 207350 92020 207650 92090
rect 207850 92020 208000 92090
rect 196000 91980 208000 92020
rect 196000 91910 196150 91980
rect 196350 91910 196650 91980
rect 196850 91910 197150 91980
rect 197350 91910 197650 91980
rect 197850 91910 198150 91980
rect 198350 91910 198650 91980
rect 198850 91910 199150 91980
rect 199350 91910 199650 91980
rect 199850 91910 200150 91980
rect 200350 91910 200650 91980
rect 200850 91910 201150 91980
rect 201350 91910 201650 91980
rect 201850 91910 202150 91980
rect 202350 91910 202650 91980
rect 202850 91910 203150 91980
rect 203350 91910 203650 91980
rect 203850 91910 204150 91980
rect 204350 91910 204650 91980
rect 204850 91910 205150 91980
rect 205350 91910 205650 91980
rect 205850 91910 206150 91980
rect 206350 91910 206650 91980
rect 206850 91910 207150 91980
rect 207350 91910 207650 91980
rect 207850 91910 208000 91980
rect 196000 91900 208000 91910
rect 196000 91880 196120 91900
rect 196380 91880 196620 91900
rect 196880 91880 197120 91900
rect 197380 91880 197620 91900
rect 197880 91880 198120 91900
rect 198380 91880 198620 91900
rect 198880 91880 199120 91900
rect 199380 91880 199620 91900
rect 199880 91880 200120 91900
rect 200380 91880 200620 91900
rect 200880 91880 201120 91900
rect 201380 91880 201620 91900
rect 201880 91880 202120 91900
rect 202380 91880 202620 91900
rect 202880 91880 203120 91900
rect 203380 91880 203620 91900
rect 203880 91880 204120 91900
rect 204380 91880 204620 91900
rect 204880 91880 205120 91900
rect 205380 91880 205620 91900
rect 205880 91880 206120 91900
rect 206380 91880 206620 91900
rect 206880 91880 207120 91900
rect 207380 91880 207620 91900
rect 207880 91880 208000 91900
rect 196000 91850 196100 91880
rect 196000 91650 196020 91850
rect 196090 91650 196100 91850
rect 196000 91620 196100 91650
rect 196400 91850 196600 91880
rect 196400 91650 196410 91850
rect 196480 91650 196520 91850
rect 196590 91650 196600 91850
rect 196400 91620 196600 91650
rect 196900 91850 197100 91880
rect 196900 91650 196910 91850
rect 196980 91650 197020 91850
rect 197090 91650 197100 91850
rect 196900 91620 197100 91650
rect 197400 91850 197600 91880
rect 197400 91650 197410 91850
rect 197480 91650 197520 91850
rect 197590 91650 197600 91850
rect 197400 91620 197600 91650
rect 197900 91850 198100 91880
rect 197900 91650 197910 91850
rect 197980 91650 198020 91850
rect 198090 91650 198100 91850
rect 197900 91620 198100 91650
rect 198400 91850 198600 91880
rect 198400 91650 198410 91850
rect 198480 91650 198520 91850
rect 198590 91650 198600 91850
rect 198400 91620 198600 91650
rect 198900 91850 199100 91880
rect 198900 91650 198910 91850
rect 198980 91650 199020 91850
rect 199090 91650 199100 91850
rect 198900 91620 199100 91650
rect 199400 91850 199600 91880
rect 199400 91650 199410 91850
rect 199480 91650 199520 91850
rect 199590 91650 199600 91850
rect 199400 91620 199600 91650
rect 199900 91850 200100 91880
rect 199900 91650 199910 91850
rect 199980 91650 200020 91850
rect 200090 91650 200100 91850
rect 199900 91620 200100 91650
rect 200400 91850 200600 91880
rect 200400 91650 200410 91850
rect 200480 91650 200520 91850
rect 200590 91650 200600 91850
rect 200400 91620 200600 91650
rect 200900 91850 201100 91880
rect 200900 91650 200910 91850
rect 200980 91650 201020 91850
rect 201090 91650 201100 91850
rect 200900 91620 201100 91650
rect 201400 91850 201600 91880
rect 201400 91650 201410 91850
rect 201480 91650 201520 91850
rect 201590 91650 201600 91850
rect 201400 91620 201600 91650
rect 201900 91850 202100 91880
rect 201900 91650 201910 91850
rect 201980 91650 202020 91850
rect 202090 91650 202100 91850
rect 201900 91620 202100 91650
rect 202400 91850 202600 91880
rect 202400 91650 202410 91850
rect 202480 91650 202520 91850
rect 202590 91650 202600 91850
rect 202400 91620 202600 91650
rect 202900 91850 203100 91880
rect 202900 91650 202910 91850
rect 202980 91650 203020 91850
rect 203090 91650 203100 91850
rect 202900 91620 203100 91650
rect 203400 91850 203600 91880
rect 203400 91650 203410 91850
rect 203480 91650 203520 91850
rect 203590 91650 203600 91850
rect 203400 91620 203600 91650
rect 203900 91850 204100 91880
rect 203900 91650 203910 91850
rect 203980 91650 204020 91850
rect 204090 91650 204100 91850
rect 203900 91620 204100 91650
rect 204400 91850 204600 91880
rect 204400 91650 204410 91850
rect 204480 91650 204520 91850
rect 204590 91650 204600 91850
rect 204400 91620 204600 91650
rect 204900 91850 205100 91880
rect 204900 91650 204910 91850
rect 204980 91650 205020 91850
rect 205090 91650 205100 91850
rect 204900 91620 205100 91650
rect 205400 91850 205600 91880
rect 205400 91650 205410 91850
rect 205480 91650 205520 91850
rect 205590 91650 205600 91850
rect 205400 91620 205600 91650
rect 205900 91850 206100 91880
rect 205900 91650 205910 91850
rect 205980 91650 206020 91850
rect 206090 91650 206100 91850
rect 205900 91620 206100 91650
rect 206400 91850 206600 91880
rect 206400 91650 206410 91850
rect 206480 91650 206520 91850
rect 206590 91650 206600 91850
rect 206400 91620 206600 91650
rect 206900 91850 207100 91880
rect 206900 91650 206910 91850
rect 206980 91650 207020 91850
rect 207090 91650 207100 91850
rect 206900 91620 207100 91650
rect 207400 91850 207600 91880
rect 207400 91650 207410 91850
rect 207480 91650 207520 91850
rect 207590 91650 207600 91850
rect 207400 91620 207600 91650
rect 207900 91850 208000 91880
rect 207900 91650 207910 91850
rect 207980 91650 208000 91850
rect 207900 91620 208000 91650
rect 196000 91600 196120 91620
rect 196380 91600 196620 91620
rect 196880 91600 197120 91620
rect 197380 91600 197620 91620
rect 197880 91600 198120 91620
rect 198380 91600 198620 91620
rect 198880 91600 199120 91620
rect 199380 91600 199620 91620
rect 199880 91600 200120 91620
rect 200380 91600 200620 91620
rect 200880 91600 201120 91620
rect 201380 91600 201620 91620
rect 201880 91600 202120 91620
rect 202380 91600 202620 91620
rect 202880 91600 203120 91620
rect 203380 91600 203620 91620
rect 203880 91600 204120 91620
rect 204380 91600 204620 91620
rect 204880 91600 205120 91620
rect 205380 91600 205620 91620
rect 205880 91600 206120 91620
rect 206380 91600 206620 91620
rect 206880 91600 207120 91620
rect 207380 91600 207620 91620
rect 207880 91600 208000 91620
rect 196000 91590 208000 91600
rect 196000 91520 196150 91590
rect 196350 91520 196650 91590
rect 196850 91520 197150 91590
rect 197350 91520 197650 91590
rect 197850 91520 198150 91590
rect 198350 91520 198650 91590
rect 198850 91520 199150 91590
rect 199350 91520 199650 91590
rect 199850 91520 200150 91590
rect 200350 91520 200650 91590
rect 200850 91520 201150 91590
rect 201350 91520 201650 91590
rect 201850 91520 202150 91590
rect 202350 91520 202650 91590
rect 202850 91520 203150 91590
rect 203350 91520 203650 91590
rect 203850 91520 204150 91590
rect 204350 91520 204650 91590
rect 204850 91520 205150 91590
rect 205350 91520 205650 91590
rect 205850 91520 206150 91590
rect 206350 91520 206650 91590
rect 206850 91520 207150 91590
rect 207350 91520 207650 91590
rect 207850 91520 208000 91590
rect 196000 91480 208000 91520
rect 196000 91410 196150 91480
rect 196350 91410 196650 91480
rect 196850 91410 197150 91480
rect 197350 91410 197650 91480
rect 197850 91410 198150 91480
rect 198350 91410 198650 91480
rect 198850 91410 199150 91480
rect 199350 91410 199650 91480
rect 199850 91410 200150 91480
rect 200350 91410 200650 91480
rect 200850 91410 201150 91480
rect 201350 91410 201650 91480
rect 201850 91410 202150 91480
rect 202350 91410 202650 91480
rect 202850 91410 203150 91480
rect 203350 91410 203650 91480
rect 203850 91410 204150 91480
rect 204350 91410 204650 91480
rect 204850 91410 205150 91480
rect 205350 91410 205650 91480
rect 205850 91410 206150 91480
rect 206350 91410 206650 91480
rect 206850 91410 207150 91480
rect 207350 91410 207650 91480
rect 207850 91410 208000 91480
rect 196000 91400 208000 91410
rect 196000 91380 196120 91400
rect 196380 91380 196620 91400
rect 196880 91380 197120 91400
rect 197380 91380 197620 91400
rect 197880 91380 198120 91400
rect 198380 91380 198620 91400
rect 198880 91380 199120 91400
rect 199380 91380 199620 91400
rect 199880 91380 200120 91400
rect 200380 91380 200620 91400
rect 200880 91380 201120 91400
rect 201380 91380 201620 91400
rect 201880 91380 202120 91400
rect 202380 91380 202620 91400
rect 202880 91380 203120 91400
rect 203380 91380 203620 91400
rect 203880 91380 204120 91400
rect 204380 91380 204620 91400
rect 204880 91380 205120 91400
rect 205380 91380 205620 91400
rect 205880 91380 206120 91400
rect 206380 91380 206620 91400
rect 206880 91380 207120 91400
rect 207380 91380 207620 91400
rect 207880 91380 208000 91400
rect 196000 91350 196100 91380
rect 196000 91150 196020 91350
rect 196090 91150 196100 91350
rect 196000 91120 196100 91150
rect 196400 91350 196600 91380
rect 196400 91150 196410 91350
rect 196480 91150 196520 91350
rect 196590 91150 196600 91350
rect 196400 91120 196600 91150
rect 196900 91350 197100 91380
rect 196900 91150 196910 91350
rect 196980 91150 197020 91350
rect 197090 91150 197100 91350
rect 196900 91120 197100 91150
rect 197400 91350 197600 91380
rect 197400 91150 197410 91350
rect 197480 91150 197520 91350
rect 197590 91150 197600 91350
rect 197400 91120 197600 91150
rect 197900 91350 198100 91380
rect 197900 91150 197910 91350
rect 197980 91150 198020 91350
rect 198090 91150 198100 91350
rect 197900 91120 198100 91150
rect 198400 91350 198600 91380
rect 198400 91150 198410 91350
rect 198480 91150 198520 91350
rect 198590 91150 198600 91350
rect 198400 91120 198600 91150
rect 198900 91350 199100 91380
rect 198900 91150 198910 91350
rect 198980 91150 199020 91350
rect 199090 91150 199100 91350
rect 198900 91120 199100 91150
rect 199400 91350 199600 91380
rect 199400 91150 199410 91350
rect 199480 91150 199520 91350
rect 199590 91150 199600 91350
rect 199400 91120 199600 91150
rect 199900 91350 200100 91380
rect 199900 91150 199910 91350
rect 199980 91150 200020 91350
rect 200090 91150 200100 91350
rect 199900 91120 200100 91150
rect 200400 91350 200600 91380
rect 200400 91150 200410 91350
rect 200480 91150 200520 91350
rect 200590 91150 200600 91350
rect 200400 91120 200600 91150
rect 200900 91350 201100 91380
rect 200900 91150 200910 91350
rect 200980 91150 201020 91350
rect 201090 91150 201100 91350
rect 200900 91120 201100 91150
rect 201400 91350 201600 91380
rect 201400 91150 201410 91350
rect 201480 91150 201520 91350
rect 201590 91150 201600 91350
rect 201400 91120 201600 91150
rect 201900 91350 202100 91380
rect 201900 91150 201910 91350
rect 201980 91150 202020 91350
rect 202090 91150 202100 91350
rect 201900 91120 202100 91150
rect 202400 91350 202600 91380
rect 202400 91150 202410 91350
rect 202480 91150 202520 91350
rect 202590 91150 202600 91350
rect 202400 91120 202600 91150
rect 202900 91350 203100 91380
rect 202900 91150 202910 91350
rect 202980 91150 203020 91350
rect 203090 91150 203100 91350
rect 202900 91120 203100 91150
rect 203400 91350 203600 91380
rect 203400 91150 203410 91350
rect 203480 91150 203520 91350
rect 203590 91150 203600 91350
rect 203400 91120 203600 91150
rect 203900 91350 204100 91380
rect 203900 91150 203910 91350
rect 203980 91150 204020 91350
rect 204090 91150 204100 91350
rect 203900 91120 204100 91150
rect 204400 91350 204600 91380
rect 204400 91150 204410 91350
rect 204480 91150 204520 91350
rect 204590 91150 204600 91350
rect 204400 91120 204600 91150
rect 204900 91350 205100 91380
rect 204900 91150 204910 91350
rect 204980 91150 205020 91350
rect 205090 91150 205100 91350
rect 204900 91120 205100 91150
rect 205400 91350 205600 91380
rect 205400 91150 205410 91350
rect 205480 91150 205520 91350
rect 205590 91150 205600 91350
rect 205400 91120 205600 91150
rect 205900 91350 206100 91380
rect 205900 91150 205910 91350
rect 205980 91150 206020 91350
rect 206090 91150 206100 91350
rect 205900 91120 206100 91150
rect 206400 91350 206600 91380
rect 206400 91150 206410 91350
rect 206480 91150 206520 91350
rect 206590 91150 206600 91350
rect 206400 91120 206600 91150
rect 206900 91350 207100 91380
rect 206900 91150 206910 91350
rect 206980 91150 207020 91350
rect 207090 91150 207100 91350
rect 206900 91120 207100 91150
rect 207400 91350 207600 91380
rect 207400 91150 207410 91350
rect 207480 91150 207520 91350
rect 207590 91150 207600 91350
rect 207400 91120 207600 91150
rect 207900 91350 208000 91380
rect 207900 91150 207910 91350
rect 207980 91150 208000 91350
rect 207900 91120 208000 91150
rect 196000 91100 196120 91120
rect 196380 91100 196620 91120
rect 196880 91100 197120 91120
rect 197380 91100 197620 91120
rect 197880 91100 198120 91120
rect 198380 91100 198620 91120
rect 198880 91100 199120 91120
rect 199380 91100 199620 91120
rect 199880 91100 200120 91120
rect 200380 91100 200620 91120
rect 200880 91100 201120 91120
rect 201380 91100 201620 91120
rect 201880 91100 202120 91120
rect 202380 91100 202620 91120
rect 202880 91100 203120 91120
rect 203380 91100 203620 91120
rect 203880 91100 204120 91120
rect 204380 91100 204620 91120
rect 204880 91100 205120 91120
rect 205380 91100 205620 91120
rect 205880 91100 206120 91120
rect 206380 91100 206620 91120
rect 206880 91100 207120 91120
rect 207380 91100 207620 91120
rect 207880 91100 208000 91120
rect 196000 91090 208000 91100
rect 196000 91020 196150 91090
rect 196350 91020 196650 91090
rect 196850 91020 197150 91090
rect 197350 91020 197650 91090
rect 197850 91020 198150 91090
rect 198350 91020 198650 91090
rect 198850 91020 199150 91090
rect 199350 91020 199650 91090
rect 199850 91020 200150 91090
rect 200350 91020 200650 91090
rect 200850 91020 201150 91090
rect 201350 91020 201650 91090
rect 201850 91020 202150 91090
rect 202350 91020 202650 91090
rect 202850 91020 203150 91090
rect 203350 91020 203650 91090
rect 203850 91020 204150 91090
rect 204350 91020 204650 91090
rect 204850 91020 205150 91090
rect 205350 91020 205650 91090
rect 205850 91020 206150 91090
rect 206350 91020 206650 91090
rect 206850 91020 207150 91090
rect 207350 91020 207650 91090
rect 207850 91020 208000 91090
rect 196000 90980 208000 91020
rect 196000 90910 196150 90980
rect 196350 90910 196650 90980
rect 196850 90910 197150 90980
rect 197350 90910 197650 90980
rect 197850 90910 198150 90980
rect 198350 90910 198650 90980
rect 198850 90910 199150 90980
rect 199350 90910 199650 90980
rect 199850 90910 200150 90980
rect 200350 90910 200650 90980
rect 200850 90910 201150 90980
rect 201350 90910 201650 90980
rect 201850 90910 202150 90980
rect 202350 90910 202650 90980
rect 202850 90910 203150 90980
rect 203350 90910 203650 90980
rect 203850 90910 204150 90980
rect 204350 90910 204650 90980
rect 204850 90910 205150 90980
rect 205350 90910 205650 90980
rect 205850 90910 206150 90980
rect 206350 90910 206650 90980
rect 206850 90910 207150 90980
rect 207350 90910 207650 90980
rect 207850 90910 208000 90980
rect 196000 90900 208000 90910
rect 196000 90880 196120 90900
rect 196380 90880 196620 90900
rect 196880 90880 197120 90900
rect 197380 90880 197620 90900
rect 197880 90880 198120 90900
rect 198380 90880 198620 90900
rect 198880 90880 199120 90900
rect 199380 90880 199620 90900
rect 199880 90880 200120 90900
rect 200380 90880 200620 90900
rect 200880 90880 201120 90900
rect 201380 90880 201620 90900
rect 201880 90880 202120 90900
rect 202380 90880 202620 90900
rect 202880 90880 203120 90900
rect 203380 90880 203620 90900
rect 203880 90880 204120 90900
rect 204380 90880 204620 90900
rect 204880 90880 205120 90900
rect 205380 90880 205620 90900
rect 205880 90880 206120 90900
rect 206380 90880 206620 90900
rect 206880 90880 207120 90900
rect 207380 90880 207620 90900
rect 207880 90880 208000 90900
rect 196000 90850 196100 90880
rect 196000 90650 196020 90850
rect 196090 90650 196100 90850
rect 196000 90620 196100 90650
rect 196400 90850 196600 90880
rect 196400 90650 196410 90850
rect 196480 90650 196520 90850
rect 196590 90650 196600 90850
rect 196400 90620 196600 90650
rect 196900 90850 197100 90880
rect 196900 90650 196910 90850
rect 196980 90650 197020 90850
rect 197090 90650 197100 90850
rect 196900 90620 197100 90650
rect 197400 90850 197600 90880
rect 197400 90650 197410 90850
rect 197480 90650 197520 90850
rect 197590 90650 197600 90850
rect 197400 90620 197600 90650
rect 197900 90850 198100 90880
rect 197900 90650 197910 90850
rect 197980 90650 198020 90850
rect 198090 90650 198100 90850
rect 197900 90620 198100 90650
rect 198400 90850 198600 90880
rect 198400 90650 198410 90850
rect 198480 90650 198520 90850
rect 198590 90650 198600 90850
rect 198400 90620 198600 90650
rect 198900 90850 199100 90880
rect 198900 90650 198910 90850
rect 198980 90650 199020 90850
rect 199090 90650 199100 90850
rect 198900 90620 199100 90650
rect 199400 90850 199600 90880
rect 199400 90650 199410 90850
rect 199480 90650 199520 90850
rect 199590 90650 199600 90850
rect 199400 90620 199600 90650
rect 199900 90850 200100 90880
rect 199900 90650 199910 90850
rect 199980 90650 200020 90850
rect 200090 90650 200100 90850
rect 199900 90620 200100 90650
rect 200400 90850 200600 90880
rect 200400 90650 200410 90850
rect 200480 90650 200520 90850
rect 200590 90650 200600 90850
rect 200400 90620 200600 90650
rect 200900 90850 201100 90880
rect 200900 90650 200910 90850
rect 200980 90650 201020 90850
rect 201090 90650 201100 90850
rect 200900 90620 201100 90650
rect 201400 90850 201600 90880
rect 201400 90650 201410 90850
rect 201480 90650 201520 90850
rect 201590 90650 201600 90850
rect 201400 90620 201600 90650
rect 201900 90850 202100 90880
rect 201900 90650 201910 90850
rect 201980 90650 202020 90850
rect 202090 90650 202100 90850
rect 201900 90620 202100 90650
rect 202400 90850 202600 90880
rect 202400 90650 202410 90850
rect 202480 90650 202520 90850
rect 202590 90650 202600 90850
rect 202400 90620 202600 90650
rect 202900 90850 203100 90880
rect 202900 90650 202910 90850
rect 202980 90650 203020 90850
rect 203090 90650 203100 90850
rect 202900 90620 203100 90650
rect 203400 90850 203600 90880
rect 203400 90650 203410 90850
rect 203480 90650 203520 90850
rect 203590 90650 203600 90850
rect 203400 90620 203600 90650
rect 203900 90850 204100 90880
rect 203900 90650 203910 90850
rect 203980 90650 204020 90850
rect 204090 90650 204100 90850
rect 203900 90620 204100 90650
rect 204400 90850 204600 90880
rect 204400 90650 204410 90850
rect 204480 90650 204520 90850
rect 204590 90650 204600 90850
rect 204400 90620 204600 90650
rect 204900 90850 205100 90880
rect 204900 90650 204910 90850
rect 204980 90650 205020 90850
rect 205090 90650 205100 90850
rect 204900 90620 205100 90650
rect 205400 90850 205600 90880
rect 205400 90650 205410 90850
rect 205480 90650 205520 90850
rect 205590 90650 205600 90850
rect 205400 90620 205600 90650
rect 205900 90850 206100 90880
rect 205900 90650 205910 90850
rect 205980 90650 206020 90850
rect 206090 90650 206100 90850
rect 205900 90620 206100 90650
rect 206400 90850 206600 90880
rect 206400 90650 206410 90850
rect 206480 90650 206520 90850
rect 206590 90650 206600 90850
rect 206400 90620 206600 90650
rect 206900 90850 207100 90880
rect 206900 90650 206910 90850
rect 206980 90650 207020 90850
rect 207090 90650 207100 90850
rect 206900 90620 207100 90650
rect 207400 90850 207600 90880
rect 207400 90650 207410 90850
rect 207480 90650 207520 90850
rect 207590 90650 207600 90850
rect 207400 90620 207600 90650
rect 207900 90850 208000 90880
rect 207900 90650 207910 90850
rect 207980 90650 208000 90850
rect 207900 90620 208000 90650
rect 196000 90600 196120 90620
rect 196380 90600 196620 90620
rect 196880 90600 197120 90620
rect 197380 90600 197620 90620
rect 197880 90600 198120 90620
rect 198380 90600 198620 90620
rect 198880 90600 199120 90620
rect 199380 90600 199620 90620
rect 199880 90600 200120 90620
rect 200380 90600 200620 90620
rect 200880 90600 201120 90620
rect 201380 90600 201620 90620
rect 201880 90600 202120 90620
rect 202380 90600 202620 90620
rect 202880 90600 203120 90620
rect 203380 90600 203620 90620
rect 203880 90600 204120 90620
rect 204380 90600 204620 90620
rect 204880 90600 205120 90620
rect 205380 90600 205620 90620
rect 205880 90600 206120 90620
rect 206380 90600 206620 90620
rect 206880 90600 207120 90620
rect 207380 90600 207620 90620
rect 207880 90600 208000 90620
rect 196000 90590 208000 90600
rect 196000 90520 196150 90590
rect 196350 90520 196650 90590
rect 196850 90520 197150 90590
rect 197350 90520 197650 90590
rect 197850 90520 198150 90590
rect 198350 90520 198650 90590
rect 198850 90520 199150 90590
rect 199350 90520 199650 90590
rect 199850 90520 200150 90590
rect 200350 90520 200650 90590
rect 200850 90520 201150 90590
rect 201350 90520 201650 90590
rect 201850 90520 202150 90590
rect 202350 90520 202650 90590
rect 202850 90520 203150 90590
rect 203350 90520 203650 90590
rect 203850 90520 204150 90590
rect 204350 90520 204650 90590
rect 204850 90520 205150 90590
rect 205350 90520 205650 90590
rect 205850 90520 206150 90590
rect 206350 90520 206650 90590
rect 206850 90520 207150 90590
rect 207350 90520 207650 90590
rect 207850 90520 208000 90590
rect 196000 90480 208000 90520
rect 196000 90410 196150 90480
rect 196350 90410 196650 90480
rect 196850 90410 197150 90480
rect 197350 90410 197650 90480
rect 197850 90410 198150 90480
rect 198350 90410 198650 90480
rect 198850 90410 199150 90480
rect 199350 90410 199650 90480
rect 199850 90410 200150 90480
rect 200350 90410 200650 90480
rect 200850 90410 201150 90480
rect 201350 90410 201650 90480
rect 201850 90410 202150 90480
rect 202350 90410 202650 90480
rect 202850 90410 203150 90480
rect 203350 90410 203650 90480
rect 203850 90410 204150 90480
rect 204350 90410 204650 90480
rect 204850 90410 205150 90480
rect 205350 90410 205650 90480
rect 205850 90410 206150 90480
rect 206350 90410 206650 90480
rect 206850 90410 207150 90480
rect 207350 90410 207650 90480
rect 207850 90410 208000 90480
rect 196000 90400 208000 90410
rect 196000 90380 196120 90400
rect 196380 90380 196620 90400
rect 196880 90380 197120 90400
rect 197380 90380 197620 90400
rect 197880 90380 198120 90400
rect 198380 90380 198620 90400
rect 198880 90380 199120 90400
rect 199380 90380 199620 90400
rect 199880 90380 200120 90400
rect 200380 90380 200620 90400
rect 200880 90380 201120 90400
rect 201380 90380 201620 90400
rect 201880 90380 202120 90400
rect 202380 90380 202620 90400
rect 202880 90380 203120 90400
rect 203380 90380 203620 90400
rect 203880 90380 204120 90400
rect 204380 90380 204620 90400
rect 204880 90380 205120 90400
rect 205380 90380 205620 90400
rect 205880 90380 206120 90400
rect 206380 90380 206620 90400
rect 206880 90380 207120 90400
rect 207380 90380 207620 90400
rect 207880 90380 208000 90400
rect 196000 90350 196100 90380
rect 196000 90150 196020 90350
rect 196090 90150 196100 90350
rect 196000 90120 196100 90150
rect 196400 90350 196600 90380
rect 196400 90150 196410 90350
rect 196480 90150 196520 90350
rect 196590 90150 196600 90350
rect 196400 90120 196600 90150
rect 196900 90350 197100 90380
rect 196900 90150 196910 90350
rect 196980 90150 197020 90350
rect 197090 90150 197100 90350
rect 196900 90120 197100 90150
rect 197400 90350 197600 90380
rect 197400 90150 197410 90350
rect 197480 90150 197520 90350
rect 197590 90150 197600 90350
rect 197400 90120 197600 90150
rect 197900 90350 198100 90380
rect 197900 90150 197910 90350
rect 197980 90150 198020 90350
rect 198090 90150 198100 90350
rect 197900 90120 198100 90150
rect 198400 90350 198600 90380
rect 198400 90150 198410 90350
rect 198480 90150 198520 90350
rect 198590 90150 198600 90350
rect 198400 90120 198600 90150
rect 198900 90350 199100 90380
rect 198900 90150 198910 90350
rect 198980 90150 199020 90350
rect 199090 90150 199100 90350
rect 198900 90120 199100 90150
rect 199400 90350 199600 90380
rect 199400 90150 199410 90350
rect 199480 90150 199520 90350
rect 199590 90150 199600 90350
rect 199400 90120 199600 90150
rect 199900 90350 200100 90380
rect 199900 90150 199910 90350
rect 199980 90150 200020 90350
rect 200090 90150 200100 90350
rect 199900 90120 200100 90150
rect 200400 90350 200600 90380
rect 200400 90150 200410 90350
rect 200480 90150 200520 90350
rect 200590 90150 200600 90350
rect 200400 90120 200600 90150
rect 200900 90350 201100 90380
rect 200900 90150 200910 90350
rect 200980 90150 201020 90350
rect 201090 90150 201100 90350
rect 200900 90120 201100 90150
rect 201400 90350 201600 90380
rect 201400 90150 201410 90350
rect 201480 90150 201520 90350
rect 201590 90150 201600 90350
rect 201400 90120 201600 90150
rect 201900 90350 202100 90380
rect 201900 90150 201910 90350
rect 201980 90150 202020 90350
rect 202090 90150 202100 90350
rect 201900 90120 202100 90150
rect 202400 90350 202600 90380
rect 202400 90150 202410 90350
rect 202480 90150 202520 90350
rect 202590 90150 202600 90350
rect 202400 90120 202600 90150
rect 202900 90350 203100 90380
rect 202900 90150 202910 90350
rect 202980 90150 203020 90350
rect 203090 90150 203100 90350
rect 202900 90120 203100 90150
rect 203400 90350 203600 90380
rect 203400 90150 203410 90350
rect 203480 90150 203520 90350
rect 203590 90150 203600 90350
rect 203400 90120 203600 90150
rect 203900 90350 204100 90380
rect 203900 90150 203910 90350
rect 203980 90150 204020 90350
rect 204090 90150 204100 90350
rect 203900 90120 204100 90150
rect 204400 90350 204600 90380
rect 204400 90150 204410 90350
rect 204480 90150 204520 90350
rect 204590 90150 204600 90350
rect 204400 90120 204600 90150
rect 204900 90350 205100 90380
rect 204900 90150 204910 90350
rect 204980 90150 205020 90350
rect 205090 90150 205100 90350
rect 204900 90120 205100 90150
rect 205400 90350 205600 90380
rect 205400 90150 205410 90350
rect 205480 90150 205520 90350
rect 205590 90150 205600 90350
rect 205400 90120 205600 90150
rect 205900 90350 206100 90380
rect 205900 90150 205910 90350
rect 205980 90150 206020 90350
rect 206090 90150 206100 90350
rect 205900 90120 206100 90150
rect 206400 90350 206600 90380
rect 206400 90150 206410 90350
rect 206480 90150 206520 90350
rect 206590 90150 206600 90350
rect 206400 90120 206600 90150
rect 206900 90350 207100 90380
rect 206900 90150 206910 90350
rect 206980 90150 207020 90350
rect 207090 90150 207100 90350
rect 206900 90120 207100 90150
rect 207400 90350 207600 90380
rect 207400 90150 207410 90350
rect 207480 90150 207520 90350
rect 207590 90150 207600 90350
rect 207400 90120 207600 90150
rect 207900 90350 208000 90380
rect 207900 90150 207910 90350
rect 207980 90150 208000 90350
rect 207900 90120 208000 90150
rect 196000 90100 196120 90120
rect 196380 90100 196620 90120
rect 196880 90100 197120 90120
rect 197380 90100 197620 90120
rect 197880 90100 198120 90120
rect 198380 90100 198620 90120
rect 198880 90100 199120 90120
rect 199380 90100 199620 90120
rect 199880 90100 200120 90120
rect 200380 90100 200620 90120
rect 200880 90100 201120 90120
rect 201380 90100 201620 90120
rect 201880 90100 202120 90120
rect 202380 90100 202620 90120
rect 202880 90100 203120 90120
rect 203380 90100 203620 90120
rect 203880 90100 204120 90120
rect 204380 90100 204620 90120
rect 204880 90100 205120 90120
rect 205380 90100 205620 90120
rect 205880 90100 206120 90120
rect 206380 90100 206620 90120
rect 206880 90100 207120 90120
rect 207380 90100 207620 90120
rect 207880 90100 208000 90120
rect 196000 90090 208000 90100
rect 196000 90020 196150 90090
rect 196350 90020 196650 90090
rect 196850 90020 197150 90090
rect 197350 90020 197650 90090
rect 197850 90020 198150 90090
rect 198350 90020 198650 90090
rect 198850 90020 199150 90090
rect 199350 90020 199650 90090
rect 199850 90020 200150 90090
rect 200350 90020 200650 90090
rect 200850 90020 201150 90090
rect 201350 90020 201650 90090
rect 201850 90020 202150 90090
rect 202350 90020 202650 90090
rect 202850 90020 203150 90090
rect 203350 90020 203650 90090
rect 203850 90020 204150 90090
rect 204350 90020 204650 90090
rect 204850 90020 205150 90090
rect 205350 90020 205650 90090
rect 205850 90020 206150 90090
rect 206350 90020 206650 90090
rect 206850 90020 207150 90090
rect 207350 90020 207650 90090
rect 207850 90020 208000 90090
rect 196000 89980 208000 90020
rect 196000 89910 196150 89980
rect 196350 89910 196650 89980
rect 196850 89910 197150 89980
rect 197350 89910 197650 89980
rect 197850 89910 198150 89980
rect 198350 89910 198650 89980
rect 198850 89910 199150 89980
rect 199350 89910 199650 89980
rect 199850 89910 200150 89980
rect 200350 89910 200650 89980
rect 200850 89910 201150 89980
rect 201350 89910 201650 89980
rect 201850 89910 202150 89980
rect 202350 89910 202650 89980
rect 202850 89910 203150 89980
rect 203350 89910 203650 89980
rect 203850 89910 204150 89980
rect 204350 89910 204650 89980
rect 204850 89910 205150 89980
rect 205350 89910 205650 89980
rect 205850 89910 206150 89980
rect 206350 89910 206650 89980
rect 206850 89910 207150 89980
rect 207350 89910 207650 89980
rect 207850 89910 208000 89980
rect 196000 89900 208000 89910
rect 196000 89880 196120 89900
rect 196380 89880 196620 89900
rect 196880 89880 197120 89900
rect 197380 89880 197620 89900
rect 197880 89880 198120 89900
rect 198380 89880 198620 89900
rect 198880 89880 199120 89900
rect 199380 89880 199620 89900
rect 199880 89880 200120 89900
rect 200380 89880 200620 89900
rect 200880 89880 201120 89900
rect 201380 89880 201620 89900
rect 201880 89880 202120 89900
rect 202380 89880 202620 89900
rect 202880 89880 203120 89900
rect 203380 89880 203620 89900
rect 203880 89880 204120 89900
rect 204380 89880 204620 89900
rect 204880 89880 205120 89900
rect 205380 89880 205620 89900
rect 205880 89880 206120 89900
rect 206380 89880 206620 89900
rect 206880 89880 207120 89900
rect 207380 89880 207620 89900
rect 207880 89880 208000 89900
rect 196000 89850 196100 89880
rect 196000 89650 196020 89850
rect 196090 89650 196100 89850
rect 196000 89620 196100 89650
rect 196400 89850 196600 89880
rect 196400 89650 196410 89850
rect 196480 89650 196520 89850
rect 196590 89650 196600 89850
rect 196400 89620 196600 89650
rect 196900 89850 197100 89880
rect 196900 89650 196910 89850
rect 196980 89650 197020 89850
rect 197090 89650 197100 89850
rect 196900 89620 197100 89650
rect 197400 89850 197600 89880
rect 197400 89650 197410 89850
rect 197480 89650 197520 89850
rect 197590 89650 197600 89850
rect 197400 89620 197600 89650
rect 197900 89850 198100 89880
rect 197900 89650 197910 89850
rect 197980 89650 198020 89850
rect 198090 89650 198100 89850
rect 197900 89620 198100 89650
rect 198400 89850 198600 89880
rect 198400 89650 198410 89850
rect 198480 89650 198520 89850
rect 198590 89650 198600 89850
rect 198400 89620 198600 89650
rect 198900 89850 199100 89880
rect 198900 89650 198910 89850
rect 198980 89650 199020 89850
rect 199090 89650 199100 89850
rect 198900 89620 199100 89650
rect 199400 89850 199600 89880
rect 199400 89650 199410 89850
rect 199480 89650 199520 89850
rect 199590 89650 199600 89850
rect 199400 89620 199600 89650
rect 199900 89850 200100 89880
rect 199900 89650 199910 89850
rect 199980 89650 200020 89850
rect 200090 89650 200100 89850
rect 199900 89620 200100 89650
rect 200400 89850 200600 89880
rect 200400 89650 200410 89850
rect 200480 89650 200520 89850
rect 200590 89650 200600 89850
rect 200400 89620 200600 89650
rect 200900 89850 201100 89880
rect 200900 89650 200910 89850
rect 200980 89650 201020 89850
rect 201090 89650 201100 89850
rect 200900 89620 201100 89650
rect 201400 89850 201600 89880
rect 201400 89650 201410 89850
rect 201480 89650 201520 89850
rect 201590 89650 201600 89850
rect 201400 89620 201600 89650
rect 201900 89850 202100 89880
rect 201900 89650 201910 89850
rect 201980 89650 202020 89850
rect 202090 89650 202100 89850
rect 201900 89620 202100 89650
rect 202400 89850 202600 89880
rect 202400 89650 202410 89850
rect 202480 89650 202520 89850
rect 202590 89650 202600 89850
rect 202400 89620 202600 89650
rect 202900 89850 203100 89880
rect 202900 89650 202910 89850
rect 202980 89650 203020 89850
rect 203090 89650 203100 89850
rect 202900 89620 203100 89650
rect 203400 89850 203600 89880
rect 203400 89650 203410 89850
rect 203480 89650 203520 89850
rect 203590 89650 203600 89850
rect 203400 89620 203600 89650
rect 203900 89850 204100 89880
rect 203900 89650 203910 89850
rect 203980 89650 204020 89850
rect 204090 89650 204100 89850
rect 203900 89620 204100 89650
rect 204400 89850 204600 89880
rect 204400 89650 204410 89850
rect 204480 89650 204520 89850
rect 204590 89650 204600 89850
rect 204400 89620 204600 89650
rect 204900 89850 205100 89880
rect 204900 89650 204910 89850
rect 204980 89650 205020 89850
rect 205090 89650 205100 89850
rect 204900 89620 205100 89650
rect 205400 89850 205600 89880
rect 205400 89650 205410 89850
rect 205480 89650 205520 89850
rect 205590 89650 205600 89850
rect 205400 89620 205600 89650
rect 205900 89850 206100 89880
rect 205900 89650 205910 89850
rect 205980 89650 206020 89850
rect 206090 89650 206100 89850
rect 205900 89620 206100 89650
rect 206400 89850 206600 89880
rect 206400 89650 206410 89850
rect 206480 89650 206520 89850
rect 206590 89650 206600 89850
rect 206400 89620 206600 89650
rect 206900 89850 207100 89880
rect 206900 89650 206910 89850
rect 206980 89650 207020 89850
rect 207090 89650 207100 89850
rect 206900 89620 207100 89650
rect 207400 89850 207600 89880
rect 207400 89650 207410 89850
rect 207480 89650 207520 89850
rect 207590 89650 207600 89850
rect 207400 89620 207600 89650
rect 207900 89850 208000 89880
rect 207900 89650 207910 89850
rect 207980 89650 208000 89850
rect 207900 89620 208000 89650
rect 196000 89600 196120 89620
rect 196380 89600 196620 89620
rect 196880 89600 197120 89620
rect 197380 89600 197620 89620
rect 197880 89600 198120 89620
rect 198380 89600 198620 89620
rect 198880 89600 199120 89620
rect 199380 89600 199620 89620
rect 199880 89600 200120 89620
rect 200380 89600 200620 89620
rect 200880 89600 201120 89620
rect 201380 89600 201620 89620
rect 201880 89600 202120 89620
rect 202380 89600 202620 89620
rect 202880 89600 203120 89620
rect 203380 89600 203620 89620
rect 203880 89600 204120 89620
rect 204380 89600 204620 89620
rect 204880 89600 205120 89620
rect 205380 89600 205620 89620
rect 205880 89600 206120 89620
rect 206380 89600 206620 89620
rect 206880 89600 207120 89620
rect 207380 89600 207620 89620
rect 207880 89600 208000 89620
rect 196000 89590 208000 89600
rect 196000 89520 196150 89590
rect 196350 89520 196650 89590
rect 196850 89520 197150 89590
rect 197350 89520 197650 89590
rect 197850 89520 198150 89590
rect 198350 89520 198650 89590
rect 198850 89520 199150 89590
rect 199350 89520 199650 89590
rect 199850 89520 200150 89590
rect 200350 89520 200650 89590
rect 200850 89520 201150 89590
rect 201350 89520 201650 89590
rect 201850 89520 202150 89590
rect 202350 89520 202650 89590
rect 202850 89520 203150 89590
rect 203350 89520 203650 89590
rect 203850 89520 204150 89590
rect 204350 89520 204650 89590
rect 204850 89520 205150 89590
rect 205350 89520 205650 89590
rect 205850 89520 206150 89590
rect 206350 89520 206650 89590
rect 206850 89520 207150 89590
rect 207350 89520 207650 89590
rect 207850 89520 208000 89590
rect 196000 89480 208000 89520
rect 196000 89410 196150 89480
rect 196350 89410 196650 89480
rect 196850 89410 197150 89480
rect 197350 89410 197650 89480
rect 197850 89410 198150 89480
rect 198350 89410 198650 89480
rect 198850 89410 199150 89480
rect 199350 89410 199650 89480
rect 199850 89410 200150 89480
rect 200350 89410 200650 89480
rect 200850 89410 201150 89480
rect 201350 89410 201650 89480
rect 201850 89410 202150 89480
rect 202350 89410 202650 89480
rect 202850 89410 203150 89480
rect 203350 89410 203650 89480
rect 203850 89410 204150 89480
rect 204350 89410 204650 89480
rect 204850 89410 205150 89480
rect 205350 89410 205650 89480
rect 205850 89410 206150 89480
rect 206350 89410 206650 89480
rect 206850 89410 207150 89480
rect 207350 89410 207650 89480
rect 207850 89410 208000 89480
rect 196000 89400 208000 89410
rect 196000 89380 196120 89400
rect 196380 89380 196620 89400
rect 196880 89380 197120 89400
rect 197380 89380 197620 89400
rect 197880 89380 198120 89400
rect 198380 89380 198620 89400
rect 198880 89380 199120 89400
rect 199380 89380 199620 89400
rect 199880 89380 200120 89400
rect 200380 89380 200620 89400
rect 200880 89380 201120 89400
rect 201380 89380 201620 89400
rect 201880 89380 202120 89400
rect 202380 89380 202620 89400
rect 202880 89380 203120 89400
rect 203380 89380 203620 89400
rect 203880 89380 204120 89400
rect 204380 89380 204620 89400
rect 204880 89380 205120 89400
rect 205380 89380 205620 89400
rect 205880 89380 206120 89400
rect 206380 89380 206620 89400
rect 206880 89380 207120 89400
rect 207380 89380 207620 89400
rect 207880 89380 208000 89400
rect 196000 89350 196100 89380
rect 196000 89150 196020 89350
rect 196090 89150 196100 89350
rect 196000 89120 196100 89150
rect 196400 89350 196600 89380
rect 196400 89150 196410 89350
rect 196480 89150 196520 89350
rect 196590 89150 196600 89350
rect 196400 89120 196600 89150
rect 196900 89350 197100 89380
rect 196900 89150 196910 89350
rect 196980 89150 197020 89350
rect 197090 89150 197100 89350
rect 196900 89120 197100 89150
rect 197400 89350 197600 89380
rect 197400 89150 197410 89350
rect 197480 89150 197520 89350
rect 197590 89150 197600 89350
rect 197400 89120 197600 89150
rect 197900 89350 198100 89380
rect 197900 89150 197910 89350
rect 197980 89150 198020 89350
rect 198090 89150 198100 89350
rect 197900 89120 198100 89150
rect 198400 89350 198600 89380
rect 198400 89150 198410 89350
rect 198480 89150 198520 89350
rect 198590 89150 198600 89350
rect 198400 89120 198600 89150
rect 198900 89350 199100 89380
rect 198900 89150 198910 89350
rect 198980 89150 199020 89350
rect 199090 89150 199100 89350
rect 198900 89120 199100 89150
rect 199400 89350 199600 89380
rect 199400 89150 199410 89350
rect 199480 89150 199520 89350
rect 199590 89150 199600 89350
rect 199400 89120 199600 89150
rect 199900 89350 200100 89380
rect 199900 89150 199910 89350
rect 199980 89150 200020 89350
rect 200090 89150 200100 89350
rect 199900 89120 200100 89150
rect 200400 89350 200600 89380
rect 200400 89150 200410 89350
rect 200480 89150 200520 89350
rect 200590 89150 200600 89350
rect 200400 89120 200600 89150
rect 200900 89350 201100 89380
rect 200900 89150 200910 89350
rect 200980 89150 201020 89350
rect 201090 89150 201100 89350
rect 200900 89120 201100 89150
rect 201400 89350 201600 89380
rect 201400 89150 201410 89350
rect 201480 89150 201520 89350
rect 201590 89150 201600 89350
rect 201400 89120 201600 89150
rect 201900 89350 202100 89380
rect 201900 89150 201910 89350
rect 201980 89150 202020 89350
rect 202090 89150 202100 89350
rect 201900 89120 202100 89150
rect 202400 89350 202600 89380
rect 202400 89150 202410 89350
rect 202480 89150 202520 89350
rect 202590 89150 202600 89350
rect 202400 89120 202600 89150
rect 202900 89350 203100 89380
rect 202900 89150 202910 89350
rect 202980 89150 203020 89350
rect 203090 89150 203100 89350
rect 202900 89120 203100 89150
rect 203400 89350 203600 89380
rect 203400 89150 203410 89350
rect 203480 89150 203520 89350
rect 203590 89150 203600 89350
rect 203400 89120 203600 89150
rect 203900 89350 204100 89380
rect 203900 89150 203910 89350
rect 203980 89150 204020 89350
rect 204090 89150 204100 89350
rect 203900 89120 204100 89150
rect 204400 89350 204600 89380
rect 204400 89150 204410 89350
rect 204480 89150 204520 89350
rect 204590 89150 204600 89350
rect 204400 89120 204600 89150
rect 204900 89350 205100 89380
rect 204900 89150 204910 89350
rect 204980 89150 205020 89350
rect 205090 89150 205100 89350
rect 204900 89120 205100 89150
rect 205400 89350 205600 89380
rect 205400 89150 205410 89350
rect 205480 89150 205520 89350
rect 205590 89150 205600 89350
rect 205400 89120 205600 89150
rect 205900 89350 206100 89380
rect 205900 89150 205910 89350
rect 205980 89150 206020 89350
rect 206090 89150 206100 89350
rect 205900 89120 206100 89150
rect 206400 89350 206600 89380
rect 206400 89150 206410 89350
rect 206480 89150 206520 89350
rect 206590 89150 206600 89350
rect 206400 89120 206600 89150
rect 206900 89350 207100 89380
rect 206900 89150 206910 89350
rect 206980 89150 207020 89350
rect 207090 89150 207100 89350
rect 206900 89120 207100 89150
rect 207400 89350 207600 89380
rect 207400 89150 207410 89350
rect 207480 89150 207520 89350
rect 207590 89150 207600 89350
rect 207400 89120 207600 89150
rect 207900 89350 208000 89380
rect 207900 89150 207910 89350
rect 207980 89150 208000 89350
rect 207900 89120 208000 89150
rect 196000 89100 196120 89120
rect 196380 89100 196620 89120
rect 196880 89100 197120 89120
rect 197380 89100 197620 89120
rect 197880 89100 198120 89120
rect 198380 89100 198620 89120
rect 198880 89100 199120 89120
rect 199380 89100 199620 89120
rect 199880 89100 200120 89120
rect 200380 89100 200620 89120
rect 200880 89100 201120 89120
rect 201380 89100 201620 89120
rect 201880 89100 202120 89120
rect 202380 89100 202620 89120
rect 202880 89100 203120 89120
rect 203380 89100 203620 89120
rect 203880 89100 204120 89120
rect 204380 89100 204620 89120
rect 204880 89100 205120 89120
rect 205380 89100 205620 89120
rect 205880 89100 206120 89120
rect 206380 89100 206620 89120
rect 206880 89100 207120 89120
rect 207380 89100 207620 89120
rect 207880 89100 208000 89120
rect 196000 89090 208000 89100
rect 196000 89020 196150 89090
rect 196350 89020 196650 89090
rect 196850 89020 197150 89090
rect 197350 89020 197650 89090
rect 197850 89020 198150 89090
rect 198350 89020 198650 89090
rect 198850 89020 199150 89090
rect 199350 89020 199650 89090
rect 199850 89020 200150 89090
rect 200350 89020 200650 89090
rect 200850 89020 201150 89090
rect 201350 89020 201650 89090
rect 201850 89020 202150 89090
rect 202350 89020 202650 89090
rect 202850 89020 203150 89090
rect 203350 89020 203650 89090
rect 203850 89020 204150 89090
rect 204350 89020 204650 89090
rect 204850 89020 205150 89090
rect 205350 89020 205650 89090
rect 205850 89020 206150 89090
rect 206350 89020 206650 89090
rect 206850 89020 207150 89090
rect 207350 89020 207650 89090
rect 207850 89020 208000 89090
rect 196000 88980 208000 89020
rect 196000 88910 196150 88980
rect 196350 88910 196650 88980
rect 196850 88910 197150 88980
rect 197350 88910 197650 88980
rect 197850 88910 198150 88980
rect 198350 88910 198650 88980
rect 198850 88910 199150 88980
rect 199350 88910 199650 88980
rect 199850 88910 200150 88980
rect 200350 88910 200650 88980
rect 200850 88910 201150 88980
rect 201350 88910 201650 88980
rect 201850 88910 202150 88980
rect 202350 88910 202650 88980
rect 202850 88910 203150 88980
rect 203350 88910 203650 88980
rect 203850 88910 204150 88980
rect 204350 88910 204650 88980
rect 204850 88910 205150 88980
rect 205350 88910 205650 88980
rect 205850 88910 206150 88980
rect 206350 88910 206650 88980
rect 206850 88910 207150 88980
rect 207350 88910 207650 88980
rect 207850 88910 208000 88980
rect 196000 88900 208000 88910
rect 196000 88880 196120 88900
rect 196380 88880 196620 88900
rect 196880 88880 197120 88900
rect 197380 88880 197620 88900
rect 197880 88880 198120 88900
rect 198380 88880 198620 88900
rect 198880 88880 199120 88900
rect 199380 88880 199620 88900
rect 199880 88880 200120 88900
rect 200380 88880 200620 88900
rect 200880 88880 201120 88900
rect 201380 88880 201620 88900
rect 201880 88880 202120 88900
rect 202380 88880 202620 88900
rect 202880 88880 203120 88900
rect 203380 88880 203620 88900
rect 203880 88880 204120 88900
rect 204380 88880 204620 88900
rect 204880 88880 205120 88900
rect 205380 88880 205620 88900
rect 205880 88880 206120 88900
rect 206380 88880 206620 88900
rect 206880 88880 207120 88900
rect 207380 88880 207620 88900
rect 207880 88880 208000 88900
rect 196000 88850 196100 88880
rect 196000 88650 196020 88850
rect 196090 88650 196100 88850
rect 196000 88620 196100 88650
rect 196400 88850 196600 88880
rect 196400 88650 196410 88850
rect 196480 88650 196520 88850
rect 196590 88650 196600 88850
rect 196400 88620 196600 88650
rect 196900 88850 197100 88880
rect 196900 88650 196910 88850
rect 196980 88650 197020 88850
rect 197090 88650 197100 88850
rect 196900 88620 197100 88650
rect 197400 88850 197600 88880
rect 197400 88650 197410 88850
rect 197480 88650 197520 88850
rect 197590 88650 197600 88850
rect 197400 88620 197600 88650
rect 197900 88850 198100 88880
rect 197900 88650 197910 88850
rect 197980 88650 198020 88850
rect 198090 88650 198100 88850
rect 197900 88620 198100 88650
rect 198400 88850 198600 88880
rect 198400 88650 198410 88850
rect 198480 88650 198520 88850
rect 198590 88650 198600 88850
rect 198400 88620 198600 88650
rect 198900 88850 199100 88880
rect 198900 88650 198910 88850
rect 198980 88650 199020 88850
rect 199090 88650 199100 88850
rect 198900 88620 199100 88650
rect 199400 88850 199600 88880
rect 199400 88650 199410 88850
rect 199480 88650 199520 88850
rect 199590 88650 199600 88850
rect 199400 88620 199600 88650
rect 199900 88850 200100 88880
rect 199900 88650 199910 88850
rect 199980 88650 200020 88850
rect 200090 88650 200100 88850
rect 199900 88620 200100 88650
rect 200400 88850 200600 88880
rect 200400 88650 200410 88850
rect 200480 88650 200520 88850
rect 200590 88650 200600 88850
rect 200400 88620 200600 88650
rect 200900 88850 201100 88880
rect 200900 88650 200910 88850
rect 200980 88650 201020 88850
rect 201090 88650 201100 88850
rect 200900 88620 201100 88650
rect 201400 88850 201600 88880
rect 201400 88650 201410 88850
rect 201480 88650 201520 88850
rect 201590 88650 201600 88850
rect 201400 88620 201600 88650
rect 201900 88850 202100 88880
rect 201900 88650 201910 88850
rect 201980 88650 202020 88850
rect 202090 88650 202100 88850
rect 201900 88620 202100 88650
rect 202400 88850 202600 88880
rect 202400 88650 202410 88850
rect 202480 88650 202520 88850
rect 202590 88650 202600 88850
rect 202400 88620 202600 88650
rect 202900 88850 203100 88880
rect 202900 88650 202910 88850
rect 202980 88650 203020 88850
rect 203090 88650 203100 88850
rect 202900 88620 203100 88650
rect 203400 88850 203600 88880
rect 203400 88650 203410 88850
rect 203480 88650 203520 88850
rect 203590 88650 203600 88850
rect 203400 88620 203600 88650
rect 203900 88850 204100 88880
rect 203900 88650 203910 88850
rect 203980 88650 204020 88850
rect 204090 88650 204100 88850
rect 203900 88620 204100 88650
rect 204400 88850 204600 88880
rect 204400 88650 204410 88850
rect 204480 88650 204520 88850
rect 204590 88650 204600 88850
rect 204400 88620 204600 88650
rect 204900 88850 205100 88880
rect 204900 88650 204910 88850
rect 204980 88650 205020 88850
rect 205090 88650 205100 88850
rect 204900 88620 205100 88650
rect 205400 88850 205600 88880
rect 205400 88650 205410 88850
rect 205480 88650 205520 88850
rect 205590 88650 205600 88850
rect 205400 88620 205600 88650
rect 205900 88850 206100 88880
rect 205900 88650 205910 88850
rect 205980 88650 206020 88850
rect 206090 88650 206100 88850
rect 205900 88620 206100 88650
rect 206400 88850 206600 88880
rect 206400 88650 206410 88850
rect 206480 88650 206520 88850
rect 206590 88650 206600 88850
rect 206400 88620 206600 88650
rect 206900 88850 207100 88880
rect 206900 88650 206910 88850
rect 206980 88650 207020 88850
rect 207090 88650 207100 88850
rect 206900 88620 207100 88650
rect 207400 88850 207600 88880
rect 207400 88650 207410 88850
rect 207480 88650 207520 88850
rect 207590 88650 207600 88850
rect 207400 88620 207600 88650
rect 207900 88850 208000 88880
rect 207900 88650 207910 88850
rect 207980 88650 208000 88850
rect 207900 88620 208000 88650
rect 196000 88600 196120 88620
rect 196380 88600 196620 88620
rect 196880 88600 197120 88620
rect 197380 88600 197620 88620
rect 197880 88600 198120 88620
rect 198380 88600 198620 88620
rect 198880 88600 199120 88620
rect 199380 88600 199620 88620
rect 199880 88600 200120 88620
rect 200380 88600 200620 88620
rect 200880 88600 201120 88620
rect 201380 88600 201620 88620
rect 201880 88600 202120 88620
rect 202380 88600 202620 88620
rect 202880 88600 203120 88620
rect 203380 88600 203620 88620
rect 203880 88600 204120 88620
rect 204380 88600 204620 88620
rect 204880 88600 205120 88620
rect 205380 88600 205620 88620
rect 205880 88600 206120 88620
rect 206380 88600 206620 88620
rect 206880 88600 207120 88620
rect 207380 88600 207620 88620
rect 207880 88600 208000 88620
rect 196000 88590 208000 88600
rect 196000 88520 196150 88590
rect 196350 88520 196650 88590
rect 196850 88520 197150 88590
rect 197350 88520 197650 88590
rect 197850 88520 198150 88590
rect 198350 88520 198650 88590
rect 198850 88520 199150 88590
rect 199350 88520 199650 88590
rect 199850 88520 200150 88590
rect 200350 88520 200650 88590
rect 200850 88520 201150 88590
rect 201350 88520 201650 88590
rect 201850 88520 202150 88590
rect 202350 88520 202650 88590
rect 202850 88520 203150 88590
rect 203350 88520 203650 88590
rect 203850 88520 204150 88590
rect 204350 88520 204650 88590
rect 204850 88520 205150 88590
rect 205350 88520 205650 88590
rect 205850 88520 206150 88590
rect 206350 88520 206650 88590
rect 206850 88520 207150 88590
rect 207350 88520 207650 88590
rect 207850 88520 208000 88590
rect 196000 88480 208000 88520
rect 196000 88410 196150 88480
rect 196350 88410 196650 88480
rect 196850 88410 197150 88480
rect 197350 88410 197650 88480
rect 197850 88410 198150 88480
rect 198350 88410 198650 88480
rect 198850 88410 199150 88480
rect 199350 88410 199650 88480
rect 199850 88410 200150 88480
rect 200350 88410 200650 88480
rect 200850 88410 201150 88480
rect 201350 88410 201650 88480
rect 201850 88410 202150 88480
rect 202350 88410 202650 88480
rect 202850 88410 203150 88480
rect 203350 88410 203650 88480
rect 203850 88410 204150 88480
rect 204350 88410 204650 88480
rect 204850 88410 205150 88480
rect 205350 88410 205650 88480
rect 205850 88410 206150 88480
rect 206350 88410 206650 88480
rect 206850 88410 207150 88480
rect 207350 88410 207650 88480
rect 207850 88410 208000 88480
rect 196000 88400 208000 88410
rect 196000 88380 196120 88400
rect 196380 88380 196620 88400
rect 196880 88380 197120 88400
rect 197380 88380 197620 88400
rect 197880 88380 198120 88400
rect 198380 88380 198620 88400
rect 198880 88380 199120 88400
rect 199380 88380 199620 88400
rect 199880 88380 200120 88400
rect 200380 88380 200620 88400
rect 200880 88380 201120 88400
rect 201380 88380 201620 88400
rect 201880 88380 202120 88400
rect 202380 88380 202620 88400
rect 202880 88380 203120 88400
rect 203380 88380 203620 88400
rect 203880 88380 204120 88400
rect 204380 88380 204620 88400
rect 204880 88380 205120 88400
rect 205380 88380 205620 88400
rect 205880 88380 206120 88400
rect 206380 88380 206620 88400
rect 206880 88380 207120 88400
rect 207380 88380 207620 88400
rect 207880 88380 208000 88400
rect 196000 88350 196100 88380
rect 196000 88150 196020 88350
rect 196090 88150 196100 88350
rect 196000 88120 196100 88150
rect 196400 88350 196600 88380
rect 196400 88150 196410 88350
rect 196480 88150 196520 88350
rect 196590 88150 196600 88350
rect 196400 88120 196600 88150
rect 196900 88350 197100 88380
rect 196900 88150 196910 88350
rect 196980 88150 197020 88350
rect 197090 88150 197100 88350
rect 196900 88120 197100 88150
rect 197400 88350 197600 88380
rect 197400 88150 197410 88350
rect 197480 88150 197520 88350
rect 197590 88150 197600 88350
rect 197400 88120 197600 88150
rect 197900 88350 198100 88380
rect 197900 88150 197910 88350
rect 197980 88150 198020 88350
rect 198090 88150 198100 88350
rect 197900 88120 198100 88150
rect 198400 88350 198600 88380
rect 198400 88150 198410 88350
rect 198480 88150 198520 88350
rect 198590 88150 198600 88350
rect 198400 88120 198600 88150
rect 198900 88350 199100 88380
rect 198900 88150 198910 88350
rect 198980 88150 199020 88350
rect 199090 88150 199100 88350
rect 198900 88120 199100 88150
rect 199400 88350 199600 88380
rect 199400 88150 199410 88350
rect 199480 88150 199520 88350
rect 199590 88150 199600 88350
rect 199400 88120 199600 88150
rect 199900 88350 200100 88380
rect 199900 88150 199910 88350
rect 199980 88150 200020 88350
rect 200090 88150 200100 88350
rect 199900 88120 200100 88150
rect 200400 88350 200600 88380
rect 200400 88150 200410 88350
rect 200480 88150 200520 88350
rect 200590 88150 200600 88350
rect 200400 88120 200600 88150
rect 200900 88350 201100 88380
rect 200900 88150 200910 88350
rect 200980 88150 201020 88350
rect 201090 88150 201100 88350
rect 200900 88120 201100 88150
rect 201400 88350 201600 88380
rect 201400 88150 201410 88350
rect 201480 88150 201520 88350
rect 201590 88150 201600 88350
rect 201400 88120 201600 88150
rect 201900 88350 202100 88380
rect 201900 88150 201910 88350
rect 201980 88150 202020 88350
rect 202090 88150 202100 88350
rect 201900 88120 202100 88150
rect 202400 88350 202600 88380
rect 202400 88150 202410 88350
rect 202480 88150 202520 88350
rect 202590 88150 202600 88350
rect 202400 88120 202600 88150
rect 202900 88350 203100 88380
rect 202900 88150 202910 88350
rect 202980 88150 203020 88350
rect 203090 88150 203100 88350
rect 202900 88120 203100 88150
rect 203400 88350 203600 88380
rect 203400 88150 203410 88350
rect 203480 88150 203520 88350
rect 203590 88150 203600 88350
rect 203400 88120 203600 88150
rect 203900 88350 204100 88380
rect 203900 88150 203910 88350
rect 203980 88150 204020 88350
rect 204090 88150 204100 88350
rect 203900 88120 204100 88150
rect 204400 88350 204600 88380
rect 204400 88150 204410 88350
rect 204480 88150 204520 88350
rect 204590 88150 204600 88350
rect 204400 88120 204600 88150
rect 204900 88350 205100 88380
rect 204900 88150 204910 88350
rect 204980 88150 205020 88350
rect 205090 88150 205100 88350
rect 204900 88120 205100 88150
rect 205400 88350 205600 88380
rect 205400 88150 205410 88350
rect 205480 88150 205520 88350
rect 205590 88150 205600 88350
rect 205400 88120 205600 88150
rect 205900 88350 206100 88380
rect 205900 88150 205910 88350
rect 205980 88150 206020 88350
rect 206090 88150 206100 88350
rect 205900 88120 206100 88150
rect 206400 88350 206600 88380
rect 206400 88150 206410 88350
rect 206480 88150 206520 88350
rect 206590 88150 206600 88350
rect 206400 88120 206600 88150
rect 206900 88350 207100 88380
rect 206900 88150 206910 88350
rect 206980 88150 207020 88350
rect 207090 88150 207100 88350
rect 206900 88120 207100 88150
rect 207400 88350 207600 88380
rect 207400 88150 207410 88350
rect 207480 88150 207520 88350
rect 207590 88150 207600 88350
rect 207400 88120 207600 88150
rect 207900 88350 208000 88380
rect 207900 88150 207910 88350
rect 207980 88150 208000 88350
rect 207900 88120 208000 88150
rect 196000 88100 196120 88120
rect 196380 88100 196620 88120
rect 196880 88100 197120 88120
rect 197380 88100 197620 88120
rect 197880 88100 198120 88120
rect 198380 88100 198620 88120
rect 198880 88100 199120 88120
rect 199380 88100 199620 88120
rect 199880 88100 200120 88120
rect 200380 88100 200620 88120
rect 200880 88100 201120 88120
rect 201380 88100 201620 88120
rect 201880 88100 202120 88120
rect 202380 88100 202620 88120
rect 202880 88100 203120 88120
rect 203380 88100 203620 88120
rect 203880 88100 204120 88120
rect 204380 88100 204620 88120
rect 204880 88100 205120 88120
rect 205380 88100 205620 88120
rect 205880 88100 206120 88120
rect 206380 88100 206620 88120
rect 206880 88100 207120 88120
rect 207380 88100 207620 88120
rect 207880 88100 208000 88120
rect 196000 88090 208000 88100
rect 196000 88020 196150 88090
rect 196350 88020 196650 88090
rect 196850 88020 197150 88090
rect 197350 88020 197650 88090
rect 197850 88020 198150 88090
rect 198350 88020 198650 88090
rect 198850 88020 199150 88090
rect 199350 88020 199650 88090
rect 199850 88020 200150 88090
rect 200350 88020 200650 88090
rect 200850 88020 201150 88090
rect 201350 88020 201650 88090
rect 201850 88020 202150 88090
rect 202350 88020 202650 88090
rect 202850 88020 203150 88090
rect 203350 88020 203650 88090
rect 203850 88020 204150 88090
rect 204350 88020 204650 88090
rect 204850 88020 205150 88090
rect 205350 88020 205650 88090
rect 205850 88020 206150 88090
rect 206350 88020 206650 88090
rect 206850 88020 207150 88090
rect 207350 88020 207650 88090
rect 207850 88020 208000 88090
rect 196000 87980 208000 88020
rect 196000 87910 196150 87980
rect 196350 87910 196650 87980
rect 196850 87910 197150 87980
rect 197350 87910 197650 87980
rect 197850 87910 198150 87980
rect 198350 87910 198650 87980
rect 198850 87910 199150 87980
rect 199350 87910 199650 87980
rect 199850 87910 200150 87980
rect 200350 87910 200650 87980
rect 200850 87910 201150 87980
rect 201350 87910 201650 87980
rect 201850 87910 202150 87980
rect 202350 87910 202650 87980
rect 202850 87910 203150 87980
rect 203350 87910 203650 87980
rect 203850 87910 204150 87980
rect 204350 87910 204650 87980
rect 204850 87910 205150 87980
rect 205350 87910 205650 87980
rect 205850 87910 206150 87980
rect 206350 87910 206650 87980
rect 206850 87910 207150 87980
rect 207350 87910 207650 87980
rect 207850 87910 208000 87980
rect 196000 87900 208000 87910
rect 196000 87880 196120 87900
rect 196380 87880 196620 87900
rect 196880 87880 197120 87900
rect 197380 87880 197620 87900
rect 197880 87880 198120 87900
rect 198380 87880 198620 87900
rect 198880 87880 199120 87900
rect 199380 87880 199620 87900
rect 199880 87880 200120 87900
rect 200380 87880 200620 87900
rect 200880 87880 201120 87900
rect 201380 87880 201620 87900
rect 201880 87880 202120 87900
rect 202380 87880 202620 87900
rect 202880 87880 203120 87900
rect 203380 87880 203620 87900
rect 203880 87880 204120 87900
rect 204380 87880 204620 87900
rect 204880 87880 205120 87900
rect 205380 87880 205620 87900
rect 205880 87880 206120 87900
rect 206380 87880 206620 87900
rect 206880 87880 207120 87900
rect 207380 87880 207620 87900
rect 207880 87880 208000 87900
rect 196000 87850 196100 87880
rect 196000 87650 196020 87850
rect 196090 87650 196100 87850
rect 196000 87620 196100 87650
rect 196400 87850 196600 87880
rect 196400 87650 196410 87850
rect 196480 87650 196520 87850
rect 196590 87650 196600 87850
rect 196400 87620 196600 87650
rect 196900 87850 197100 87880
rect 196900 87650 196910 87850
rect 196980 87650 197020 87850
rect 197090 87650 197100 87850
rect 196900 87620 197100 87650
rect 197400 87850 197600 87880
rect 197400 87650 197410 87850
rect 197480 87650 197520 87850
rect 197590 87650 197600 87850
rect 197400 87620 197600 87650
rect 197900 87850 198100 87880
rect 197900 87650 197910 87850
rect 197980 87650 198020 87850
rect 198090 87650 198100 87850
rect 197900 87620 198100 87650
rect 198400 87850 198600 87880
rect 198400 87650 198410 87850
rect 198480 87650 198520 87850
rect 198590 87650 198600 87850
rect 198400 87620 198600 87650
rect 198900 87850 199100 87880
rect 198900 87650 198910 87850
rect 198980 87650 199020 87850
rect 199090 87650 199100 87850
rect 198900 87620 199100 87650
rect 199400 87850 199600 87880
rect 199400 87650 199410 87850
rect 199480 87650 199520 87850
rect 199590 87650 199600 87850
rect 199400 87620 199600 87650
rect 199900 87850 200100 87880
rect 199900 87650 199910 87850
rect 199980 87650 200020 87850
rect 200090 87650 200100 87850
rect 199900 87620 200100 87650
rect 200400 87850 200600 87880
rect 200400 87650 200410 87850
rect 200480 87650 200520 87850
rect 200590 87650 200600 87850
rect 200400 87620 200600 87650
rect 200900 87850 201100 87880
rect 200900 87650 200910 87850
rect 200980 87650 201020 87850
rect 201090 87650 201100 87850
rect 200900 87620 201100 87650
rect 201400 87850 201600 87880
rect 201400 87650 201410 87850
rect 201480 87650 201520 87850
rect 201590 87650 201600 87850
rect 201400 87620 201600 87650
rect 201900 87850 202100 87880
rect 201900 87650 201910 87850
rect 201980 87650 202020 87850
rect 202090 87650 202100 87850
rect 201900 87620 202100 87650
rect 202400 87850 202600 87880
rect 202400 87650 202410 87850
rect 202480 87650 202520 87850
rect 202590 87650 202600 87850
rect 202400 87620 202600 87650
rect 202900 87850 203100 87880
rect 202900 87650 202910 87850
rect 202980 87650 203020 87850
rect 203090 87650 203100 87850
rect 202900 87620 203100 87650
rect 203400 87850 203600 87880
rect 203400 87650 203410 87850
rect 203480 87650 203520 87850
rect 203590 87650 203600 87850
rect 203400 87620 203600 87650
rect 203900 87850 204100 87880
rect 203900 87650 203910 87850
rect 203980 87650 204020 87850
rect 204090 87650 204100 87850
rect 203900 87620 204100 87650
rect 204400 87850 204600 87880
rect 204400 87650 204410 87850
rect 204480 87650 204520 87850
rect 204590 87650 204600 87850
rect 204400 87620 204600 87650
rect 204900 87850 205100 87880
rect 204900 87650 204910 87850
rect 204980 87650 205020 87850
rect 205090 87650 205100 87850
rect 204900 87620 205100 87650
rect 205400 87850 205600 87880
rect 205400 87650 205410 87850
rect 205480 87650 205520 87850
rect 205590 87650 205600 87850
rect 205400 87620 205600 87650
rect 205900 87850 206100 87880
rect 205900 87650 205910 87850
rect 205980 87650 206020 87850
rect 206090 87650 206100 87850
rect 205900 87620 206100 87650
rect 206400 87850 206600 87880
rect 206400 87650 206410 87850
rect 206480 87650 206520 87850
rect 206590 87650 206600 87850
rect 206400 87620 206600 87650
rect 206900 87850 207100 87880
rect 206900 87650 206910 87850
rect 206980 87650 207020 87850
rect 207090 87650 207100 87850
rect 206900 87620 207100 87650
rect 207400 87850 207600 87880
rect 207400 87650 207410 87850
rect 207480 87650 207520 87850
rect 207590 87650 207600 87850
rect 207400 87620 207600 87650
rect 207900 87850 208000 87880
rect 207900 87650 207910 87850
rect 207980 87650 208000 87850
rect 207900 87620 208000 87650
rect 196000 87600 196120 87620
rect 196380 87600 196620 87620
rect 196880 87600 197120 87620
rect 197380 87600 197620 87620
rect 197880 87600 198120 87620
rect 198380 87600 198620 87620
rect 198880 87600 199120 87620
rect 199380 87600 199620 87620
rect 199880 87600 200120 87620
rect 200380 87600 200620 87620
rect 200880 87600 201120 87620
rect 201380 87600 201620 87620
rect 201880 87600 202120 87620
rect 202380 87600 202620 87620
rect 202880 87600 203120 87620
rect 203380 87600 203620 87620
rect 203880 87600 204120 87620
rect 204380 87600 204620 87620
rect 204880 87600 205120 87620
rect 205380 87600 205620 87620
rect 205880 87600 206120 87620
rect 206380 87600 206620 87620
rect 206880 87600 207120 87620
rect 207380 87600 207620 87620
rect 207880 87600 208000 87620
rect 196000 87590 208000 87600
rect 196000 87520 196150 87590
rect 196350 87520 196650 87590
rect 196850 87520 197150 87590
rect 197350 87520 197650 87590
rect 197850 87520 198150 87590
rect 198350 87520 198650 87590
rect 198850 87520 199150 87590
rect 199350 87520 199650 87590
rect 199850 87520 200150 87590
rect 200350 87520 200650 87590
rect 200850 87520 201150 87590
rect 201350 87520 201650 87590
rect 201850 87520 202150 87590
rect 202350 87520 202650 87590
rect 202850 87520 203150 87590
rect 203350 87520 203650 87590
rect 203850 87520 204150 87590
rect 204350 87520 204650 87590
rect 204850 87520 205150 87590
rect 205350 87520 205650 87590
rect 205850 87520 206150 87590
rect 206350 87520 206650 87590
rect 206850 87520 207150 87590
rect 207350 87520 207650 87590
rect 207850 87520 208000 87590
rect 196000 87480 208000 87520
rect 196000 87410 196150 87480
rect 196350 87410 196650 87480
rect 196850 87410 197150 87480
rect 197350 87410 197650 87480
rect 197850 87410 198150 87480
rect 198350 87410 198650 87480
rect 198850 87410 199150 87480
rect 199350 87410 199650 87480
rect 199850 87410 200150 87480
rect 200350 87410 200650 87480
rect 200850 87410 201150 87480
rect 201350 87410 201650 87480
rect 201850 87410 202150 87480
rect 202350 87410 202650 87480
rect 202850 87410 203150 87480
rect 203350 87410 203650 87480
rect 203850 87410 204150 87480
rect 204350 87410 204650 87480
rect 204850 87410 205150 87480
rect 205350 87410 205650 87480
rect 205850 87410 206150 87480
rect 206350 87410 206650 87480
rect 206850 87410 207150 87480
rect 207350 87410 207650 87480
rect 207850 87410 208000 87480
rect 196000 87400 208000 87410
rect 196000 87380 196120 87400
rect 196380 87380 196620 87400
rect 196880 87380 197120 87400
rect 197380 87380 197620 87400
rect 197880 87380 198120 87400
rect 198380 87380 198620 87400
rect 198880 87380 199120 87400
rect 199380 87380 199620 87400
rect 199880 87380 200120 87400
rect 200380 87380 200620 87400
rect 200880 87380 201120 87400
rect 201380 87380 201620 87400
rect 201880 87380 202120 87400
rect 202380 87380 202620 87400
rect 202880 87380 203120 87400
rect 203380 87380 203620 87400
rect 203880 87380 204120 87400
rect 204380 87380 204620 87400
rect 204880 87380 205120 87400
rect 205380 87380 205620 87400
rect 205880 87380 206120 87400
rect 206380 87380 206620 87400
rect 206880 87380 207120 87400
rect 207380 87380 207620 87400
rect 207880 87380 208000 87400
rect 196000 87350 196100 87380
rect 196000 87150 196020 87350
rect 196090 87150 196100 87350
rect 196000 87120 196100 87150
rect 196400 87350 196600 87380
rect 196400 87150 196410 87350
rect 196480 87150 196520 87350
rect 196590 87150 196600 87350
rect 196400 87120 196600 87150
rect 196900 87350 197100 87380
rect 196900 87150 196910 87350
rect 196980 87150 197020 87350
rect 197090 87150 197100 87350
rect 196900 87120 197100 87150
rect 197400 87350 197600 87380
rect 197400 87150 197410 87350
rect 197480 87150 197520 87350
rect 197590 87150 197600 87350
rect 197400 87120 197600 87150
rect 197900 87350 198100 87380
rect 197900 87150 197910 87350
rect 197980 87150 198020 87350
rect 198090 87150 198100 87350
rect 197900 87120 198100 87150
rect 198400 87350 198600 87380
rect 198400 87150 198410 87350
rect 198480 87150 198520 87350
rect 198590 87150 198600 87350
rect 198400 87120 198600 87150
rect 198900 87350 199100 87380
rect 198900 87150 198910 87350
rect 198980 87150 199020 87350
rect 199090 87150 199100 87350
rect 198900 87120 199100 87150
rect 199400 87350 199600 87380
rect 199400 87150 199410 87350
rect 199480 87150 199520 87350
rect 199590 87150 199600 87350
rect 199400 87120 199600 87150
rect 199900 87350 200100 87380
rect 199900 87150 199910 87350
rect 199980 87150 200020 87350
rect 200090 87150 200100 87350
rect 199900 87120 200100 87150
rect 200400 87350 200600 87380
rect 200400 87150 200410 87350
rect 200480 87150 200520 87350
rect 200590 87150 200600 87350
rect 200400 87120 200600 87150
rect 200900 87350 201100 87380
rect 200900 87150 200910 87350
rect 200980 87150 201020 87350
rect 201090 87150 201100 87350
rect 200900 87120 201100 87150
rect 201400 87350 201600 87380
rect 201400 87150 201410 87350
rect 201480 87150 201520 87350
rect 201590 87150 201600 87350
rect 201400 87120 201600 87150
rect 201900 87350 202100 87380
rect 201900 87150 201910 87350
rect 201980 87150 202020 87350
rect 202090 87150 202100 87350
rect 201900 87120 202100 87150
rect 202400 87350 202600 87380
rect 202400 87150 202410 87350
rect 202480 87150 202520 87350
rect 202590 87150 202600 87350
rect 202400 87120 202600 87150
rect 202900 87350 203100 87380
rect 202900 87150 202910 87350
rect 202980 87150 203020 87350
rect 203090 87150 203100 87350
rect 202900 87120 203100 87150
rect 203400 87350 203600 87380
rect 203400 87150 203410 87350
rect 203480 87150 203520 87350
rect 203590 87150 203600 87350
rect 203400 87120 203600 87150
rect 203900 87350 204100 87380
rect 203900 87150 203910 87350
rect 203980 87150 204020 87350
rect 204090 87150 204100 87350
rect 203900 87120 204100 87150
rect 204400 87350 204600 87380
rect 204400 87150 204410 87350
rect 204480 87150 204520 87350
rect 204590 87150 204600 87350
rect 204400 87120 204600 87150
rect 204900 87350 205100 87380
rect 204900 87150 204910 87350
rect 204980 87150 205020 87350
rect 205090 87150 205100 87350
rect 204900 87120 205100 87150
rect 205400 87350 205600 87380
rect 205400 87150 205410 87350
rect 205480 87150 205520 87350
rect 205590 87150 205600 87350
rect 205400 87120 205600 87150
rect 205900 87350 206100 87380
rect 205900 87150 205910 87350
rect 205980 87150 206020 87350
rect 206090 87150 206100 87350
rect 205900 87120 206100 87150
rect 206400 87350 206600 87380
rect 206400 87150 206410 87350
rect 206480 87150 206520 87350
rect 206590 87150 206600 87350
rect 206400 87120 206600 87150
rect 206900 87350 207100 87380
rect 206900 87150 206910 87350
rect 206980 87150 207020 87350
rect 207090 87150 207100 87350
rect 206900 87120 207100 87150
rect 207400 87350 207600 87380
rect 207400 87150 207410 87350
rect 207480 87150 207520 87350
rect 207590 87150 207600 87350
rect 207400 87120 207600 87150
rect 207900 87350 208000 87380
rect 207900 87150 207910 87350
rect 207980 87150 208000 87350
rect 207900 87120 208000 87150
rect 128750 87110 128910 87120
rect 128750 86870 128760 87110
rect 128900 86870 128910 87110
rect 128750 86860 128910 86870
rect 129070 87110 129230 87120
rect 129070 86870 129080 87110
rect 129220 86870 129230 87110
rect 129070 86860 129230 86870
rect 196000 87100 196120 87120
rect 196380 87100 196620 87120
rect 196880 87100 197120 87120
rect 197380 87100 197620 87120
rect 197880 87100 198120 87120
rect 198380 87100 198620 87120
rect 198880 87100 199120 87120
rect 199380 87100 199620 87120
rect 199880 87100 200120 87120
rect 200380 87100 200620 87120
rect 200880 87100 201120 87120
rect 201380 87100 201620 87120
rect 201880 87100 202120 87120
rect 202380 87100 202620 87120
rect 202880 87100 203120 87120
rect 203380 87100 203620 87120
rect 203880 87100 204120 87120
rect 204380 87100 204620 87120
rect 204880 87100 205120 87120
rect 205380 87100 205620 87120
rect 205880 87100 206120 87120
rect 206380 87100 206620 87120
rect 206880 87100 207120 87120
rect 207380 87100 207620 87120
rect 207880 87100 208000 87120
rect 196000 87090 208000 87100
rect 196000 87020 196150 87090
rect 196350 87020 196650 87090
rect 196850 87020 197150 87090
rect 197350 87020 197650 87090
rect 197850 87020 198150 87090
rect 198350 87020 198650 87090
rect 198850 87020 199150 87090
rect 199350 87020 199650 87090
rect 199850 87020 200150 87090
rect 200350 87020 200650 87090
rect 200850 87020 201150 87090
rect 201350 87020 201650 87090
rect 201850 87020 202150 87090
rect 202350 87020 202650 87090
rect 202850 87020 203150 87090
rect 203350 87020 203650 87090
rect 203850 87020 204150 87090
rect 204350 87020 204650 87090
rect 204850 87020 205150 87090
rect 205350 87020 205650 87090
rect 205850 87020 206150 87090
rect 206350 87020 206650 87090
rect 206850 87020 207150 87090
rect 207350 87020 207650 87090
rect 207850 87020 208000 87090
rect 196000 86980 208000 87020
rect 196000 86910 196150 86980
rect 196350 86910 196650 86980
rect 196850 86910 197150 86980
rect 197350 86910 197650 86980
rect 197850 86910 198150 86980
rect 198350 86910 198650 86980
rect 198850 86910 199150 86980
rect 199350 86910 199650 86980
rect 199850 86910 200150 86980
rect 200350 86910 200650 86980
rect 200850 86910 201150 86980
rect 201350 86910 201650 86980
rect 201850 86910 202150 86980
rect 202350 86910 202650 86980
rect 202850 86910 203150 86980
rect 203350 86910 203650 86980
rect 203850 86910 204150 86980
rect 204350 86910 204650 86980
rect 204850 86910 205150 86980
rect 205350 86910 205650 86980
rect 205850 86910 206150 86980
rect 206350 86910 206650 86980
rect 206850 86910 207150 86980
rect 207350 86910 207650 86980
rect 207850 86910 208000 86980
rect 196000 86900 208000 86910
rect 196000 86880 196120 86900
rect 196380 86880 196620 86900
rect 196880 86880 197120 86900
rect 197380 86880 197620 86900
rect 197880 86880 198120 86900
rect 198380 86880 198620 86900
rect 198880 86880 199120 86900
rect 199380 86880 199620 86900
rect 199880 86880 200120 86900
rect 200380 86880 200620 86900
rect 200880 86880 201120 86900
rect 201380 86880 201620 86900
rect 201880 86880 202120 86900
rect 202380 86880 202620 86900
rect 202880 86880 203120 86900
rect 203380 86880 203620 86900
rect 203880 86880 204120 86900
rect 204380 86880 204620 86900
rect 204880 86880 205120 86900
rect 205380 86880 205620 86900
rect 205880 86880 206120 86900
rect 206380 86880 206620 86900
rect 206880 86880 207120 86900
rect 207380 86880 207620 86900
rect 207880 86880 208000 86900
rect 128640 86640 128720 86720
rect 128750 86640 128830 86860
rect 128860 86630 129040 86720
rect 129070 86640 129150 86860
rect 196000 86850 196100 86880
rect 129180 86640 129260 86720
rect 196000 86650 196020 86850
rect 196090 86650 196100 86850
rect 128860 86510 128870 86630
rect 129030 86510 129040 86630
rect 128860 86500 129040 86510
rect 196000 86620 196100 86650
rect 196400 86850 196600 86880
rect 196400 86650 196410 86850
rect 196480 86650 196520 86850
rect 196590 86650 196600 86850
rect 196400 86620 196600 86650
rect 196900 86850 197100 86880
rect 196900 86650 196910 86850
rect 196980 86650 197020 86850
rect 197090 86650 197100 86850
rect 196900 86620 197100 86650
rect 197400 86850 197600 86880
rect 197400 86650 197410 86850
rect 197480 86650 197520 86850
rect 197590 86650 197600 86850
rect 197400 86620 197600 86650
rect 197900 86850 198100 86880
rect 197900 86650 197910 86850
rect 197980 86650 198020 86850
rect 198090 86650 198100 86850
rect 197900 86620 198100 86650
rect 198400 86850 198600 86880
rect 198400 86650 198410 86850
rect 198480 86650 198520 86850
rect 198590 86650 198600 86850
rect 198400 86620 198600 86650
rect 198900 86850 199100 86880
rect 198900 86650 198910 86850
rect 198980 86650 199020 86850
rect 199090 86650 199100 86850
rect 198900 86620 199100 86650
rect 199400 86850 199600 86880
rect 199400 86650 199410 86850
rect 199480 86650 199520 86850
rect 199590 86650 199600 86850
rect 199400 86620 199600 86650
rect 199900 86850 200100 86880
rect 199900 86650 199910 86850
rect 199980 86650 200020 86850
rect 200090 86650 200100 86850
rect 199900 86620 200100 86650
rect 200400 86850 200600 86880
rect 200400 86650 200410 86850
rect 200480 86650 200520 86850
rect 200590 86650 200600 86850
rect 200400 86620 200600 86650
rect 200900 86850 201100 86880
rect 200900 86650 200910 86850
rect 200980 86650 201020 86850
rect 201090 86650 201100 86850
rect 200900 86620 201100 86650
rect 201400 86850 201600 86880
rect 201400 86650 201410 86850
rect 201480 86650 201520 86850
rect 201590 86650 201600 86850
rect 201400 86620 201600 86650
rect 201900 86850 202100 86880
rect 201900 86650 201910 86850
rect 201980 86650 202020 86850
rect 202090 86650 202100 86850
rect 201900 86620 202100 86650
rect 202400 86850 202600 86880
rect 202400 86650 202410 86850
rect 202480 86650 202520 86850
rect 202590 86650 202600 86850
rect 202400 86620 202600 86650
rect 202900 86850 203100 86880
rect 202900 86650 202910 86850
rect 202980 86650 203020 86850
rect 203090 86650 203100 86850
rect 202900 86620 203100 86650
rect 203400 86850 203600 86880
rect 203400 86650 203410 86850
rect 203480 86650 203520 86850
rect 203590 86650 203600 86850
rect 203400 86620 203600 86650
rect 203900 86850 204100 86880
rect 203900 86650 203910 86850
rect 203980 86650 204020 86850
rect 204090 86650 204100 86850
rect 203900 86620 204100 86650
rect 204400 86850 204600 86880
rect 204400 86650 204410 86850
rect 204480 86650 204520 86850
rect 204590 86650 204600 86850
rect 204400 86620 204600 86650
rect 204900 86850 205100 86880
rect 204900 86650 204910 86850
rect 204980 86650 205020 86850
rect 205090 86650 205100 86850
rect 204900 86620 205100 86650
rect 205400 86850 205600 86880
rect 205400 86650 205410 86850
rect 205480 86650 205520 86850
rect 205590 86650 205600 86850
rect 205400 86620 205600 86650
rect 205900 86850 206100 86880
rect 205900 86650 205910 86850
rect 205980 86650 206020 86850
rect 206090 86650 206100 86850
rect 205900 86620 206100 86650
rect 206400 86850 206600 86880
rect 206400 86650 206410 86850
rect 206480 86650 206520 86850
rect 206590 86650 206600 86850
rect 206400 86620 206600 86650
rect 206900 86850 207100 86880
rect 206900 86650 206910 86850
rect 206980 86650 207020 86850
rect 207090 86650 207100 86850
rect 206900 86620 207100 86650
rect 207400 86850 207600 86880
rect 207400 86650 207410 86850
rect 207480 86650 207520 86850
rect 207590 86650 207600 86850
rect 207400 86620 207600 86650
rect 207900 86850 208000 86880
rect 207900 86650 207910 86850
rect 207980 86650 208000 86850
rect 207900 86620 208000 86650
rect 196000 86600 196120 86620
rect 196380 86600 196620 86620
rect 196880 86600 197120 86620
rect 197380 86600 197620 86620
rect 197880 86600 198120 86620
rect 198380 86600 198620 86620
rect 198880 86600 199120 86620
rect 199380 86600 199620 86620
rect 199880 86600 200120 86620
rect 200380 86600 200620 86620
rect 200880 86600 201120 86620
rect 201380 86600 201620 86620
rect 201880 86600 202120 86620
rect 202380 86600 202620 86620
rect 202880 86600 203120 86620
rect 203380 86600 203620 86620
rect 203880 86600 204120 86620
rect 204380 86600 204620 86620
rect 204880 86600 205120 86620
rect 205380 86600 205620 86620
rect 205880 86600 206120 86620
rect 206380 86600 206620 86620
rect 206880 86600 207120 86620
rect 207380 86600 207620 86620
rect 207880 86600 208000 86620
rect 196000 86590 208000 86600
rect 196000 86520 196150 86590
rect 196350 86520 196650 86590
rect 196850 86520 197150 86590
rect 197350 86520 197650 86590
rect 197850 86520 198150 86590
rect 198350 86520 198650 86590
rect 198850 86520 199150 86590
rect 199350 86520 199650 86590
rect 199850 86520 200150 86590
rect 200350 86520 200650 86590
rect 200850 86520 201150 86590
rect 201350 86520 201650 86590
rect 201850 86520 202150 86590
rect 202350 86520 202650 86590
rect 202850 86520 203150 86590
rect 203350 86520 203650 86590
rect 203850 86520 204150 86590
rect 204350 86520 204650 86590
rect 204850 86520 205150 86590
rect 205350 86520 205650 86590
rect 205850 86520 206150 86590
rect 206350 86520 206650 86590
rect 206850 86520 207150 86590
rect 207350 86520 207650 86590
rect 207850 86520 208000 86590
rect 196000 86480 208000 86520
rect 196000 86410 196150 86480
rect 196350 86410 196650 86480
rect 196850 86410 197150 86480
rect 197350 86410 197650 86480
rect 197850 86410 198150 86480
rect 198350 86410 198650 86480
rect 198850 86410 199150 86480
rect 199350 86410 199650 86480
rect 199850 86410 200150 86480
rect 200350 86410 200650 86480
rect 200850 86410 201150 86480
rect 201350 86410 201650 86480
rect 201850 86410 202150 86480
rect 202350 86410 202650 86480
rect 202850 86410 203150 86480
rect 203350 86410 203650 86480
rect 203850 86410 204150 86480
rect 204350 86410 204650 86480
rect 204850 86410 205150 86480
rect 205350 86410 205650 86480
rect 205850 86410 206150 86480
rect 206350 86410 206650 86480
rect 206850 86410 207150 86480
rect 207350 86410 207650 86480
rect 207850 86410 208000 86480
rect 196000 86400 208000 86410
rect 196000 86380 196120 86400
rect 196380 86380 196620 86400
rect 196880 86380 197120 86400
rect 197380 86380 197620 86400
rect 197880 86380 198120 86400
rect 198380 86380 198620 86400
rect 198880 86380 199120 86400
rect 199380 86380 199620 86400
rect 199880 86380 200120 86400
rect 200380 86380 200620 86400
rect 200880 86380 201120 86400
rect 201380 86380 201620 86400
rect 201880 86380 202120 86400
rect 202380 86380 202620 86400
rect 202880 86380 203120 86400
rect 203380 86380 203620 86400
rect 203880 86380 204120 86400
rect 204380 86380 204620 86400
rect 204880 86380 205120 86400
rect 205380 86380 205620 86400
rect 205880 86380 206120 86400
rect 206380 86380 206620 86400
rect 206880 86380 207120 86400
rect 207380 86380 207620 86400
rect 207880 86380 208000 86400
rect 196000 86350 196100 86380
rect 196000 86150 196020 86350
rect 196090 86150 196100 86350
rect 196000 86120 196100 86150
rect 196400 86350 196600 86380
rect 196400 86150 196410 86350
rect 196480 86150 196520 86350
rect 196590 86150 196600 86350
rect 196400 86120 196600 86150
rect 196900 86350 197100 86380
rect 196900 86150 196910 86350
rect 196980 86150 197020 86350
rect 197090 86150 197100 86350
rect 196900 86120 197100 86150
rect 197400 86350 197600 86380
rect 197400 86150 197410 86350
rect 197480 86150 197520 86350
rect 197590 86150 197600 86350
rect 197400 86120 197600 86150
rect 197900 86350 198100 86380
rect 197900 86150 197910 86350
rect 197980 86150 198020 86350
rect 198090 86150 198100 86350
rect 197900 86120 198100 86150
rect 198400 86350 198600 86380
rect 198400 86150 198410 86350
rect 198480 86150 198520 86350
rect 198590 86150 198600 86350
rect 198400 86120 198600 86150
rect 198900 86350 199100 86380
rect 198900 86150 198910 86350
rect 198980 86150 199020 86350
rect 199090 86150 199100 86350
rect 198900 86120 199100 86150
rect 199400 86350 199600 86380
rect 199400 86150 199410 86350
rect 199480 86150 199520 86350
rect 199590 86150 199600 86350
rect 199400 86120 199600 86150
rect 199900 86350 200100 86380
rect 199900 86150 199910 86350
rect 199980 86150 200020 86350
rect 200090 86150 200100 86350
rect 199900 86120 200100 86150
rect 200400 86350 200600 86380
rect 200400 86150 200410 86350
rect 200480 86150 200520 86350
rect 200590 86150 200600 86350
rect 200400 86120 200600 86150
rect 200900 86350 201100 86380
rect 200900 86150 200910 86350
rect 200980 86150 201020 86350
rect 201090 86150 201100 86350
rect 200900 86120 201100 86150
rect 201400 86350 201600 86380
rect 201400 86150 201410 86350
rect 201480 86150 201520 86350
rect 201590 86150 201600 86350
rect 201400 86120 201600 86150
rect 201900 86350 202100 86380
rect 201900 86150 201910 86350
rect 201980 86150 202020 86350
rect 202090 86150 202100 86350
rect 201900 86120 202100 86150
rect 202400 86350 202600 86380
rect 202400 86150 202410 86350
rect 202480 86150 202520 86350
rect 202590 86150 202600 86350
rect 202400 86120 202600 86150
rect 202900 86350 203100 86380
rect 202900 86150 202910 86350
rect 202980 86150 203020 86350
rect 203090 86150 203100 86350
rect 202900 86120 203100 86150
rect 203400 86350 203600 86380
rect 203400 86150 203410 86350
rect 203480 86150 203520 86350
rect 203590 86150 203600 86350
rect 203400 86120 203600 86150
rect 203900 86350 204100 86380
rect 203900 86150 203910 86350
rect 203980 86150 204020 86350
rect 204090 86150 204100 86350
rect 203900 86120 204100 86150
rect 204400 86350 204600 86380
rect 204400 86150 204410 86350
rect 204480 86150 204520 86350
rect 204590 86150 204600 86350
rect 204400 86120 204600 86150
rect 204900 86350 205100 86380
rect 204900 86150 204910 86350
rect 204980 86150 205020 86350
rect 205090 86150 205100 86350
rect 204900 86120 205100 86150
rect 205400 86350 205600 86380
rect 205400 86150 205410 86350
rect 205480 86150 205520 86350
rect 205590 86150 205600 86350
rect 205400 86120 205600 86150
rect 205900 86350 206100 86380
rect 205900 86150 205910 86350
rect 205980 86150 206020 86350
rect 206090 86150 206100 86350
rect 205900 86120 206100 86150
rect 206400 86350 206600 86380
rect 206400 86150 206410 86350
rect 206480 86150 206520 86350
rect 206590 86150 206600 86350
rect 206400 86120 206600 86150
rect 206900 86350 207100 86380
rect 206900 86150 206910 86350
rect 206980 86150 207020 86350
rect 207090 86150 207100 86350
rect 206900 86120 207100 86150
rect 207400 86350 207600 86380
rect 207400 86150 207410 86350
rect 207480 86150 207520 86350
rect 207590 86150 207600 86350
rect 207400 86120 207600 86150
rect 207900 86350 208000 86380
rect 207900 86150 207910 86350
rect 207980 86150 208000 86350
rect 207900 86120 208000 86150
rect 196000 86100 196120 86120
rect 196380 86100 196620 86120
rect 196880 86100 197120 86120
rect 197380 86100 197620 86120
rect 197880 86100 198120 86120
rect 198380 86100 198620 86120
rect 198880 86100 199120 86120
rect 199380 86100 199620 86120
rect 199880 86100 200120 86120
rect 200380 86100 200620 86120
rect 200880 86100 201120 86120
rect 201380 86100 201620 86120
rect 201880 86100 202120 86120
rect 202380 86100 202620 86120
rect 202880 86100 203120 86120
rect 203380 86100 203620 86120
rect 203880 86100 204120 86120
rect 204380 86100 204620 86120
rect 204880 86100 205120 86120
rect 205380 86100 205620 86120
rect 205880 86100 206120 86120
rect 206380 86100 206620 86120
rect 206880 86100 207120 86120
rect 207380 86100 207620 86120
rect 207880 86100 208000 86120
rect 196000 86090 208000 86100
rect 196000 86020 196150 86090
rect 196350 86020 196650 86090
rect 196850 86020 197150 86090
rect 197350 86020 197650 86090
rect 197850 86020 198150 86090
rect 198350 86020 198650 86090
rect 198850 86020 199150 86090
rect 199350 86020 199650 86090
rect 199850 86020 200150 86090
rect 200350 86020 200650 86090
rect 200850 86020 201150 86090
rect 201350 86020 201650 86090
rect 201850 86020 202150 86090
rect 202350 86020 202650 86090
rect 202850 86020 203150 86090
rect 203350 86020 203650 86090
rect 203850 86020 204150 86090
rect 204350 86020 204650 86090
rect 204850 86020 205150 86090
rect 205350 86020 205650 86090
rect 205850 86020 206150 86090
rect 206350 86020 206650 86090
rect 206850 86020 207150 86090
rect 207350 86020 207650 86090
rect 207850 86020 208000 86090
rect 196000 85980 208000 86020
rect 196000 85910 196150 85980
rect 196350 85910 196650 85980
rect 196850 85910 197150 85980
rect 197350 85910 197650 85980
rect 197850 85910 198150 85980
rect 198350 85910 198650 85980
rect 198850 85910 199150 85980
rect 199350 85910 199650 85980
rect 199850 85910 200150 85980
rect 200350 85910 200650 85980
rect 200850 85910 201150 85980
rect 201350 85910 201650 85980
rect 201850 85910 202150 85980
rect 202350 85910 202650 85980
rect 202850 85910 203150 85980
rect 203350 85910 203650 85980
rect 203850 85910 204150 85980
rect 204350 85910 204650 85980
rect 204850 85910 205150 85980
rect 205350 85910 205650 85980
rect 205850 85910 206150 85980
rect 206350 85910 206650 85980
rect 206850 85910 207150 85980
rect 207350 85910 207650 85980
rect 207850 85910 208000 85980
rect 196000 85900 208000 85910
rect 196000 85880 196120 85900
rect 196380 85880 196620 85900
rect 196880 85880 197120 85900
rect 197380 85880 197620 85900
rect 197880 85880 198120 85900
rect 198380 85880 198620 85900
rect 198880 85880 199120 85900
rect 199380 85880 199620 85900
rect 199880 85880 200120 85900
rect 200380 85880 200620 85900
rect 200880 85880 201120 85900
rect 201380 85880 201620 85900
rect 201880 85880 202120 85900
rect 202380 85880 202620 85900
rect 202880 85880 203120 85900
rect 203380 85880 203620 85900
rect 203880 85880 204120 85900
rect 204380 85880 204620 85900
rect 204880 85880 205120 85900
rect 205380 85880 205620 85900
rect 205880 85880 206120 85900
rect 206380 85880 206620 85900
rect 206880 85880 207120 85900
rect 207380 85880 207620 85900
rect 207880 85880 208000 85900
rect 196000 85850 196100 85880
rect 196000 85650 196020 85850
rect 196090 85650 196100 85850
rect 196000 85620 196100 85650
rect 196400 85850 196600 85880
rect 196400 85650 196410 85850
rect 196480 85650 196520 85850
rect 196590 85650 196600 85850
rect 196400 85620 196600 85650
rect 196900 85850 197100 85880
rect 196900 85650 196910 85850
rect 196980 85650 197020 85850
rect 197090 85650 197100 85850
rect 196900 85620 197100 85650
rect 197400 85850 197600 85880
rect 197400 85650 197410 85850
rect 197480 85650 197520 85850
rect 197590 85650 197600 85850
rect 197400 85620 197600 85650
rect 197900 85850 198100 85880
rect 197900 85650 197910 85850
rect 197980 85650 198020 85850
rect 198090 85650 198100 85850
rect 197900 85620 198100 85650
rect 198400 85850 198600 85880
rect 198400 85650 198410 85850
rect 198480 85650 198520 85850
rect 198590 85650 198600 85850
rect 198400 85620 198600 85650
rect 198900 85850 199100 85880
rect 198900 85650 198910 85850
rect 198980 85650 199020 85850
rect 199090 85650 199100 85850
rect 198900 85620 199100 85650
rect 199400 85850 199600 85880
rect 199400 85650 199410 85850
rect 199480 85650 199520 85850
rect 199590 85650 199600 85850
rect 199400 85620 199600 85650
rect 199900 85850 200100 85880
rect 199900 85650 199910 85850
rect 199980 85650 200020 85850
rect 200090 85650 200100 85850
rect 199900 85620 200100 85650
rect 200400 85850 200600 85880
rect 200400 85650 200410 85850
rect 200480 85650 200520 85850
rect 200590 85650 200600 85850
rect 200400 85620 200600 85650
rect 200900 85850 201100 85880
rect 200900 85650 200910 85850
rect 200980 85650 201020 85850
rect 201090 85650 201100 85850
rect 200900 85620 201100 85650
rect 201400 85850 201600 85880
rect 201400 85650 201410 85850
rect 201480 85650 201520 85850
rect 201590 85650 201600 85850
rect 201400 85620 201600 85650
rect 201900 85850 202100 85880
rect 201900 85650 201910 85850
rect 201980 85650 202020 85850
rect 202090 85650 202100 85850
rect 201900 85620 202100 85650
rect 202400 85850 202600 85880
rect 202400 85650 202410 85850
rect 202480 85650 202520 85850
rect 202590 85650 202600 85850
rect 202400 85620 202600 85650
rect 202900 85850 203100 85880
rect 202900 85650 202910 85850
rect 202980 85650 203020 85850
rect 203090 85650 203100 85850
rect 202900 85620 203100 85650
rect 203400 85850 203600 85880
rect 203400 85650 203410 85850
rect 203480 85650 203520 85850
rect 203590 85650 203600 85850
rect 203400 85620 203600 85650
rect 203900 85850 204100 85880
rect 203900 85650 203910 85850
rect 203980 85650 204020 85850
rect 204090 85650 204100 85850
rect 203900 85620 204100 85650
rect 204400 85850 204600 85880
rect 204400 85650 204410 85850
rect 204480 85650 204520 85850
rect 204590 85650 204600 85850
rect 204400 85620 204600 85650
rect 204900 85850 205100 85880
rect 204900 85650 204910 85850
rect 204980 85650 205020 85850
rect 205090 85650 205100 85850
rect 204900 85620 205100 85650
rect 205400 85850 205600 85880
rect 205400 85650 205410 85850
rect 205480 85650 205520 85850
rect 205590 85650 205600 85850
rect 205400 85620 205600 85650
rect 205900 85850 206100 85880
rect 205900 85650 205910 85850
rect 205980 85650 206020 85850
rect 206090 85650 206100 85850
rect 205900 85620 206100 85650
rect 206400 85850 206600 85880
rect 206400 85650 206410 85850
rect 206480 85650 206520 85850
rect 206590 85650 206600 85850
rect 206400 85620 206600 85650
rect 206900 85850 207100 85880
rect 206900 85650 206910 85850
rect 206980 85650 207020 85850
rect 207090 85650 207100 85850
rect 206900 85620 207100 85650
rect 207400 85850 207600 85880
rect 207400 85650 207410 85850
rect 207480 85650 207520 85850
rect 207590 85650 207600 85850
rect 207400 85620 207600 85650
rect 207900 85850 208000 85880
rect 207900 85650 207910 85850
rect 207980 85650 208000 85850
rect 207900 85620 208000 85650
rect 196000 85600 196120 85620
rect 196380 85600 196620 85620
rect 196880 85600 197120 85620
rect 197380 85600 197620 85620
rect 197880 85600 198120 85620
rect 198380 85600 198620 85620
rect 198880 85600 199120 85620
rect 199380 85600 199620 85620
rect 199880 85600 200120 85620
rect 200380 85600 200620 85620
rect 200880 85600 201120 85620
rect 201380 85600 201620 85620
rect 201880 85600 202120 85620
rect 202380 85600 202620 85620
rect 202880 85600 203120 85620
rect 203380 85600 203620 85620
rect 203880 85600 204120 85620
rect 204380 85600 204620 85620
rect 204880 85600 205120 85620
rect 205380 85600 205620 85620
rect 205880 85600 206120 85620
rect 206380 85600 206620 85620
rect 206880 85600 207120 85620
rect 207380 85600 207620 85620
rect 207880 85600 208000 85620
rect 196000 85590 208000 85600
rect 196000 85520 196150 85590
rect 196350 85520 196650 85590
rect 196850 85520 197150 85590
rect 197350 85520 197650 85590
rect 197850 85520 198150 85590
rect 198350 85520 198650 85590
rect 198850 85520 199150 85590
rect 199350 85520 199650 85590
rect 199850 85520 200150 85590
rect 200350 85520 200650 85590
rect 200850 85520 201150 85590
rect 201350 85520 201650 85590
rect 201850 85520 202150 85590
rect 202350 85520 202650 85590
rect 202850 85520 203150 85590
rect 203350 85520 203650 85590
rect 203850 85520 204150 85590
rect 204350 85520 204650 85590
rect 204850 85520 205150 85590
rect 205350 85520 205650 85590
rect 205850 85520 206150 85590
rect 206350 85520 206650 85590
rect 206850 85520 207150 85590
rect 207350 85520 207650 85590
rect 207850 85520 208000 85590
rect 196000 85480 208000 85520
rect 196000 85410 196150 85480
rect 196350 85410 196650 85480
rect 196850 85410 197150 85480
rect 197350 85410 197650 85480
rect 197850 85410 198150 85480
rect 198350 85410 198650 85480
rect 198850 85410 199150 85480
rect 199350 85410 199650 85480
rect 199850 85410 200150 85480
rect 200350 85410 200650 85480
rect 200850 85410 201150 85480
rect 201350 85410 201650 85480
rect 201850 85410 202150 85480
rect 202350 85410 202650 85480
rect 202850 85410 203150 85480
rect 203350 85410 203650 85480
rect 203850 85410 204150 85480
rect 204350 85410 204650 85480
rect 204850 85410 205150 85480
rect 205350 85410 205650 85480
rect 205850 85410 206150 85480
rect 206350 85410 206650 85480
rect 206850 85410 207150 85480
rect 207350 85410 207650 85480
rect 207850 85410 208000 85480
rect 196000 85400 208000 85410
rect 196000 85380 196120 85400
rect 196380 85380 196620 85400
rect 196880 85380 197120 85400
rect 197380 85380 197620 85400
rect 197880 85380 198120 85400
rect 198380 85380 198620 85400
rect 198880 85380 199120 85400
rect 199380 85380 199620 85400
rect 199880 85380 200120 85400
rect 200380 85380 200620 85400
rect 200880 85380 201120 85400
rect 201380 85380 201620 85400
rect 201880 85380 202120 85400
rect 202380 85380 202620 85400
rect 202880 85380 203120 85400
rect 203380 85380 203620 85400
rect 203880 85380 204120 85400
rect 204380 85380 204620 85400
rect 204880 85380 205120 85400
rect 205380 85380 205620 85400
rect 205880 85380 206120 85400
rect 206380 85380 206620 85400
rect 206880 85380 207120 85400
rect 207380 85380 207620 85400
rect 207880 85380 208000 85400
rect 196000 85350 196100 85380
rect 128640 85160 128720 85240
rect 128750 85160 128930 85240
rect 128970 85160 129150 85240
rect 129180 85160 129260 85240
rect 196000 85150 196020 85350
rect 196090 85150 196100 85350
rect 196000 85120 196100 85150
rect 196400 85350 196600 85380
rect 196400 85150 196410 85350
rect 196480 85150 196520 85350
rect 196590 85150 196600 85350
rect 196400 85120 196600 85150
rect 196900 85350 197100 85380
rect 196900 85150 196910 85350
rect 196980 85150 197020 85350
rect 197090 85150 197100 85350
rect 196900 85120 197100 85150
rect 197400 85350 197600 85380
rect 197400 85150 197410 85350
rect 197480 85150 197520 85350
rect 197590 85150 197600 85350
rect 197400 85120 197600 85150
rect 197900 85350 198100 85380
rect 197900 85150 197910 85350
rect 197980 85150 198020 85350
rect 198090 85150 198100 85350
rect 197900 85120 198100 85150
rect 198400 85350 198600 85380
rect 198400 85150 198410 85350
rect 198480 85150 198520 85350
rect 198590 85150 198600 85350
rect 198400 85120 198600 85150
rect 198900 85350 199100 85380
rect 198900 85150 198910 85350
rect 198980 85150 199020 85350
rect 199090 85150 199100 85350
rect 198900 85120 199100 85150
rect 199400 85350 199600 85380
rect 199400 85150 199410 85350
rect 199480 85150 199520 85350
rect 199590 85150 199600 85350
rect 199400 85120 199600 85150
rect 199900 85350 200100 85380
rect 199900 85150 199910 85350
rect 199980 85150 200020 85350
rect 200090 85150 200100 85350
rect 199900 85120 200100 85150
rect 200400 85350 200600 85380
rect 200400 85150 200410 85350
rect 200480 85150 200520 85350
rect 200590 85150 200600 85350
rect 200400 85120 200600 85150
rect 200900 85350 201100 85380
rect 200900 85150 200910 85350
rect 200980 85150 201020 85350
rect 201090 85150 201100 85350
rect 200900 85120 201100 85150
rect 201400 85350 201600 85380
rect 201400 85150 201410 85350
rect 201480 85150 201520 85350
rect 201590 85150 201600 85350
rect 201400 85120 201600 85150
rect 201900 85350 202100 85380
rect 201900 85150 201910 85350
rect 201980 85150 202020 85350
rect 202090 85150 202100 85350
rect 201900 85120 202100 85150
rect 202400 85350 202600 85380
rect 202400 85150 202410 85350
rect 202480 85150 202520 85350
rect 202590 85150 202600 85350
rect 202400 85120 202600 85150
rect 202900 85350 203100 85380
rect 202900 85150 202910 85350
rect 202980 85150 203020 85350
rect 203090 85150 203100 85350
rect 202900 85120 203100 85150
rect 203400 85350 203600 85380
rect 203400 85150 203410 85350
rect 203480 85150 203520 85350
rect 203590 85150 203600 85350
rect 203400 85120 203600 85150
rect 203900 85350 204100 85380
rect 203900 85150 203910 85350
rect 203980 85150 204020 85350
rect 204090 85150 204100 85350
rect 203900 85120 204100 85150
rect 204400 85350 204600 85380
rect 204400 85150 204410 85350
rect 204480 85150 204520 85350
rect 204590 85150 204600 85350
rect 204400 85120 204600 85150
rect 204900 85350 205100 85380
rect 204900 85150 204910 85350
rect 204980 85150 205020 85350
rect 205090 85150 205100 85350
rect 204900 85120 205100 85150
rect 205400 85350 205600 85380
rect 205400 85150 205410 85350
rect 205480 85150 205520 85350
rect 205590 85150 205600 85350
rect 205400 85120 205600 85150
rect 205900 85350 206100 85380
rect 205900 85150 205910 85350
rect 205980 85150 206020 85350
rect 206090 85150 206100 85350
rect 205900 85120 206100 85150
rect 206400 85350 206600 85380
rect 206400 85150 206410 85350
rect 206480 85150 206520 85350
rect 206590 85150 206600 85350
rect 206400 85120 206600 85150
rect 206900 85350 207100 85380
rect 206900 85150 206910 85350
rect 206980 85150 207020 85350
rect 207090 85150 207100 85350
rect 206900 85120 207100 85150
rect 207400 85350 207600 85380
rect 207400 85150 207410 85350
rect 207480 85150 207520 85350
rect 207590 85150 207600 85350
rect 207400 85120 207600 85150
rect 207900 85350 208000 85380
rect 207900 85150 207910 85350
rect 207980 85150 208000 85350
rect 207900 85120 208000 85150
rect 196000 85100 196120 85120
rect 196380 85100 196620 85120
rect 196880 85100 197120 85120
rect 197380 85100 197620 85120
rect 197880 85100 198120 85120
rect 198380 85100 198620 85120
rect 198880 85100 199120 85120
rect 199380 85100 199620 85120
rect 199880 85100 200120 85120
rect 200380 85100 200620 85120
rect 200880 85100 201120 85120
rect 201380 85100 201620 85120
rect 201880 85100 202120 85120
rect 202380 85100 202620 85120
rect 202880 85100 203120 85120
rect 203380 85100 203620 85120
rect 203880 85100 204120 85120
rect 204380 85100 204620 85120
rect 204880 85100 205120 85120
rect 205380 85100 205620 85120
rect 205880 85100 206120 85120
rect 206380 85100 206620 85120
rect 206880 85100 207120 85120
rect 207380 85100 207620 85120
rect 207880 85100 208000 85120
rect 196000 85090 208000 85100
rect 128520 85060 129360 85070
rect 128520 84970 128550 85060
rect 129330 84970 129360 85060
rect 196000 85020 196150 85090
rect 196350 85020 196650 85090
rect 196850 85020 197150 85090
rect 197350 85020 197650 85090
rect 197850 85020 198150 85090
rect 198350 85020 198650 85090
rect 198850 85020 199150 85090
rect 199350 85020 199650 85090
rect 199850 85020 200150 85090
rect 200350 85020 200650 85090
rect 200850 85020 201150 85090
rect 201350 85020 201650 85090
rect 201850 85020 202150 85090
rect 202350 85020 202650 85090
rect 202850 85020 203150 85090
rect 203350 85020 203650 85090
rect 203850 85020 204150 85090
rect 204350 85020 204650 85090
rect 204850 85020 205150 85090
rect 205350 85020 205650 85090
rect 205850 85020 206150 85090
rect 206350 85020 206650 85090
rect 206850 85020 207150 85090
rect 207350 85020 207650 85090
rect 207850 85020 208000 85090
rect 131120 84990 131900 85000
rect 128520 84960 129360 84970
rect 131100 84910 131910 84990
rect 196000 84980 208000 85020
rect 196000 84910 196150 84980
rect 196350 84910 196650 84980
rect 196850 84910 197150 84980
rect 197350 84910 197650 84980
rect 197850 84910 198150 84980
rect 198350 84910 198650 84980
rect 198850 84910 199150 84980
rect 199350 84910 199650 84980
rect 199850 84910 200150 84980
rect 200350 84910 200650 84980
rect 200850 84910 201150 84980
rect 201350 84910 201650 84980
rect 201850 84910 202150 84980
rect 202350 84910 202650 84980
rect 202850 84910 203150 84980
rect 203350 84910 203650 84980
rect 203850 84910 204150 84980
rect 204350 84910 204650 84980
rect 204850 84910 205150 84980
rect 205350 84910 205650 84980
rect 205850 84910 206150 84980
rect 206350 84910 206650 84980
rect 206850 84910 207150 84980
rect 207350 84910 207650 84980
rect 207850 84910 208000 84980
rect 196000 84900 208000 84910
rect 196000 84880 196120 84900
rect 196380 84880 196620 84900
rect 196880 84880 197120 84900
rect 197380 84880 197620 84900
rect 197880 84880 198120 84900
rect 198380 84880 198620 84900
rect 198880 84880 199120 84900
rect 199380 84880 199620 84900
rect 199880 84880 200120 84900
rect 200380 84880 200620 84900
rect 200880 84880 201120 84900
rect 201380 84880 201620 84900
rect 201880 84880 202120 84900
rect 202380 84880 202620 84900
rect 202880 84880 203120 84900
rect 203380 84880 203620 84900
rect 203880 84880 204120 84900
rect 204380 84880 204620 84900
rect 204880 84880 205120 84900
rect 205380 84880 205620 84900
rect 205880 84880 206120 84900
rect 206380 84880 206620 84900
rect 206880 84880 207120 84900
rect 207380 84880 207620 84900
rect 207880 84880 208000 84900
rect 196000 84850 196100 84880
rect 196000 84650 196020 84850
rect 196090 84650 196100 84850
rect 196000 84620 196100 84650
rect 196400 84850 196600 84880
rect 196400 84650 196410 84850
rect 196480 84650 196520 84850
rect 196590 84650 196600 84850
rect 196400 84620 196600 84650
rect 196900 84850 197100 84880
rect 196900 84650 196910 84850
rect 196980 84650 197020 84850
rect 197090 84650 197100 84850
rect 196900 84620 197100 84650
rect 197400 84850 197600 84880
rect 197400 84650 197410 84850
rect 197480 84650 197520 84850
rect 197590 84650 197600 84850
rect 197400 84620 197600 84650
rect 197900 84850 198100 84880
rect 197900 84650 197910 84850
rect 197980 84650 198020 84850
rect 198090 84650 198100 84850
rect 197900 84620 198100 84650
rect 198400 84850 198600 84880
rect 198400 84650 198410 84850
rect 198480 84650 198520 84850
rect 198590 84650 198600 84850
rect 198400 84620 198600 84650
rect 198900 84850 199100 84880
rect 198900 84650 198910 84850
rect 198980 84650 199020 84850
rect 199090 84650 199100 84850
rect 198900 84620 199100 84650
rect 199400 84850 199600 84880
rect 199400 84650 199410 84850
rect 199480 84650 199520 84850
rect 199590 84650 199600 84850
rect 199400 84620 199600 84650
rect 199900 84850 200100 84880
rect 199900 84650 199910 84850
rect 199980 84650 200020 84850
rect 200090 84650 200100 84850
rect 199900 84620 200100 84650
rect 200400 84850 200600 84880
rect 200400 84650 200410 84850
rect 200480 84650 200520 84850
rect 200590 84650 200600 84850
rect 200400 84620 200600 84650
rect 200900 84850 201100 84880
rect 200900 84650 200910 84850
rect 200980 84650 201020 84850
rect 201090 84650 201100 84850
rect 200900 84620 201100 84650
rect 201400 84850 201600 84880
rect 201400 84650 201410 84850
rect 201480 84650 201520 84850
rect 201590 84650 201600 84850
rect 201400 84620 201600 84650
rect 201900 84850 202100 84880
rect 201900 84650 201910 84850
rect 201980 84650 202020 84850
rect 202090 84650 202100 84850
rect 201900 84620 202100 84650
rect 202400 84850 202600 84880
rect 202400 84650 202410 84850
rect 202480 84650 202520 84850
rect 202590 84650 202600 84850
rect 202400 84620 202600 84650
rect 202900 84850 203100 84880
rect 202900 84650 202910 84850
rect 202980 84650 203020 84850
rect 203090 84650 203100 84850
rect 202900 84620 203100 84650
rect 203400 84850 203600 84880
rect 203400 84650 203410 84850
rect 203480 84650 203520 84850
rect 203590 84650 203600 84850
rect 203400 84620 203600 84650
rect 203900 84850 204100 84880
rect 203900 84650 203910 84850
rect 203980 84650 204020 84850
rect 204090 84650 204100 84850
rect 203900 84620 204100 84650
rect 204400 84850 204600 84880
rect 204400 84650 204410 84850
rect 204480 84650 204520 84850
rect 204590 84650 204600 84850
rect 204400 84620 204600 84650
rect 204900 84850 205100 84880
rect 204900 84650 204910 84850
rect 204980 84650 205020 84850
rect 205090 84650 205100 84850
rect 204900 84620 205100 84650
rect 205400 84850 205600 84880
rect 205400 84650 205410 84850
rect 205480 84650 205520 84850
rect 205590 84650 205600 84850
rect 205400 84620 205600 84650
rect 205900 84850 206100 84880
rect 205900 84650 205910 84850
rect 205980 84650 206020 84850
rect 206090 84650 206100 84850
rect 205900 84620 206100 84650
rect 206400 84850 206600 84880
rect 206400 84650 206410 84850
rect 206480 84650 206520 84850
rect 206590 84650 206600 84850
rect 206400 84620 206600 84650
rect 206900 84850 207100 84880
rect 206900 84650 206910 84850
rect 206980 84650 207020 84850
rect 207090 84650 207100 84850
rect 206900 84620 207100 84650
rect 207400 84850 207600 84880
rect 207400 84650 207410 84850
rect 207480 84650 207520 84850
rect 207590 84650 207600 84850
rect 207400 84620 207600 84650
rect 207900 84850 208000 84880
rect 207900 84650 207910 84850
rect 207980 84650 208000 84850
rect 207900 84620 208000 84650
rect 196000 84600 196120 84620
rect 196380 84600 196620 84620
rect 196880 84600 197120 84620
rect 197380 84600 197620 84620
rect 197880 84600 198120 84620
rect 198380 84600 198620 84620
rect 198880 84600 199120 84620
rect 199380 84600 199620 84620
rect 199880 84600 200120 84620
rect 200380 84600 200620 84620
rect 200880 84600 201120 84620
rect 201380 84600 201620 84620
rect 201880 84600 202120 84620
rect 202380 84600 202620 84620
rect 202880 84600 203120 84620
rect 203380 84600 203620 84620
rect 203880 84600 204120 84620
rect 204380 84600 204620 84620
rect 204880 84600 205120 84620
rect 205380 84600 205620 84620
rect 205880 84600 206120 84620
rect 206380 84600 206620 84620
rect 206880 84600 207120 84620
rect 207380 84600 207620 84620
rect 207880 84600 208000 84620
rect 196000 84590 208000 84600
rect 196000 84520 196150 84590
rect 196350 84520 196650 84590
rect 196850 84520 197150 84590
rect 197350 84520 197650 84590
rect 197850 84520 198150 84590
rect 198350 84520 198650 84590
rect 198850 84520 199150 84590
rect 199350 84520 199650 84590
rect 199850 84520 200150 84590
rect 200350 84520 200650 84590
rect 200850 84520 201150 84590
rect 201350 84520 201650 84590
rect 201850 84520 202150 84590
rect 202350 84520 202650 84590
rect 202850 84520 203150 84590
rect 203350 84520 203650 84590
rect 203850 84520 204150 84590
rect 204350 84520 204650 84590
rect 204850 84520 205150 84590
rect 205350 84520 205650 84590
rect 205850 84520 206150 84590
rect 206350 84520 206650 84590
rect 206850 84520 207150 84590
rect 207350 84520 207650 84590
rect 207850 84520 208000 84590
rect 196000 84480 208000 84520
rect 196000 84410 196150 84480
rect 196350 84410 196650 84480
rect 196850 84410 197150 84480
rect 197350 84410 197650 84480
rect 197850 84410 198150 84480
rect 198350 84410 198650 84480
rect 198850 84410 199150 84480
rect 199350 84410 199650 84480
rect 199850 84410 200150 84480
rect 200350 84410 200650 84480
rect 200850 84410 201150 84480
rect 201350 84410 201650 84480
rect 201850 84410 202150 84480
rect 202350 84410 202650 84480
rect 202850 84410 203150 84480
rect 203350 84410 203650 84480
rect 203850 84410 204150 84480
rect 204350 84410 204650 84480
rect 204850 84410 205150 84480
rect 205350 84410 205650 84480
rect 205850 84410 206150 84480
rect 206350 84410 206650 84480
rect 206850 84410 207150 84480
rect 207350 84410 207650 84480
rect 207850 84410 208000 84480
rect 196000 84400 208000 84410
rect 196000 84380 196120 84400
rect 196380 84380 196620 84400
rect 196880 84380 197120 84400
rect 197380 84380 197620 84400
rect 197880 84380 198120 84400
rect 198380 84380 198620 84400
rect 198880 84380 199120 84400
rect 199380 84380 199620 84400
rect 199880 84380 200120 84400
rect 200380 84380 200620 84400
rect 200880 84380 201120 84400
rect 201380 84380 201620 84400
rect 201880 84380 202120 84400
rect 202380 84380 202620 84400
rect 202880 84380 203120 84400
rect 203380 84380 203620 84400
rect 203880 84380 204120 84400
rect 204380 84380 204620 84400
rect 204880 84380 205120 84400
rect 205380 84380 205620 84400
rect 205880 84380 206120 84400
rect 206380 84380 206620 84400
rect 206880 84380 207120 84400
rect 207380 84380 207620 84400
rect 207880 84380 208000 84400
rect 196000 84350 196100 84380
rect 196000 84150 196020 84350
rect 196090 84150 196100 84350
rect 196000 84120 196100 84150
rect 196400 84350 196600 84380
rect 196400 84150 196410 84350
rect 196480 84150 196520 84350
rect 196590 84150 196600 84350
rect 196400 84120 196600 84150
rect 196900 84350 197100 84380
rect 196900 84150 196910 84350
rect 196980 84150 197020 84350
rect 197090 84150 197100 84350
rect 196900 84120 197100 84150
rect 197400 84350 197600 84380
rect 197400 84150 197410 84350
rect 197480 84150 197520 84350
rect 197590 84150 197600 84350
rect 197400 84120 197600 84150
rect 197900 84350 198100 84380
rect 197900 84150 197910 84350
rect 197980 84150 198020 84350
rect 198090 84150 198100 84350
rect 197900 84120 198100 84150
rect 198400 84350 198600 84380
rect 198400 84150 198410 84350
rect 198480 84150 198520 84350
rect 198590 84150 198600 84350
rect 198400 84120 198600 84150
rect 198900 84350 199100 84380
rect 198900 84150 198910 84350
rect 198980 84150 199020 84350
rect 199090 84150 199100 84350
rect 198900 84120 199100 84150
rect 199400 84350 199600 84380
rect 199400 84150 199410 84350
rect 199480 84150 199520 84350
rect 199590 84150 199600 84350
rect 199400 84120 199600 84150
rect 199900 84350 200100 84380
rect 199900 84150 199910 84350
rect 199980 84150 200020 84350
rect 200090 84150 200100 84350
rect 199900 84120 200100 84150
rect 200400 84350 200600 84380
rect 200400 84150 200410 84350
rect 200480 84150 200520 84350
rect 200590 84150 200600 84350
rect 200400 84120 200600 84150
rect 200900 84350 201100 84380
rect 200900 84150 200910 84350
rect 200980 84150 201020 84350
rect 201090 84150 201100 84350
rect 200900 84120 201100 84150
rect 201400 84350 201600 84380
rect 201400 84150 201410 84350
rect 201480 84150 201520 84350
rect 201590 84150 201600 84350
rect 201400 84120 201600 84150
rect 201900 84350 202100 84380
rect 201900 84150 201910 84350
rect 201980 84150 202020 84350
rect 202090 84150 202100 84350
rect 201900 84120 202100 84150
rect 202400 84350 202600 84380
rect 202400 84150 202410 84350
rect 202480 84150 202520 84350
rect 202590 84150 202600 84350
rect 202400 84120 202600 84150
rect 202900 84350 203100 84380
rect 202900 84150 202910 84350
rect 202980 84150 203020 84350
rect 203090 84150 203100 84350
rect 202900 84120 203100 84150
rect 203400 84350 203600 84380
rect 203400 84150 203410 84350
rect 203480 84150 203520 84350
rect 203590 84150 203600 84350
rect 203400 84120 203600 84150
rect 203900 84350 204100 84380
rect 203900 84150 203910 84350
rect 203980 84150 204020 84350
rect 204090 84150 204100 84350
rect 203900 84120 204100 84150
rect 204400 84350 204600 84380
rect 204400 84150 204410 84350
rect 204480 84150 204520 84350
rect 204590 84150 204600 84350
rect 204400 84120 204600 84150
rect 204900 84350 205100 84380
rect 204900 84150 204910 84350
rect 204980 84150 205020 84350
rect 205090 84150 205100 84350
rect 204900 84120 205100 84150
rect 205400 84350 205600 84380
rect 205400 84150 205410 84350
rect 205480 84150 205520 84350
rect 205590 84150 205600 84350
rect 205400 84120 205600 84150
rect 205900 84350 206100 84380
rect 205900 84150 205910 84350
rect 205980 84150 206020 84350
rect 206090 84150 206100 84350
rect 205900 84120 206100 84150
rect 206400 84350 206600 84380
rect 206400 84150 206410 84350
rect 206480 84150 206520 84350
rect 206590 84150 206600 84350
rect 206400 84120 206600 84150
rect 206900 84350 207100 84380
rect 206900 84150 206910 84350
rect 206980 84150 207020 84350
rect 207090 84150 207100 84350
rect 206900 84120 207100 84150
rect 207400 84350 207600 84380
rect 207400 84150 207410 84350
rect 207480 84150 207520 84350
rect 207590 84150 207600 84350
rect 207400 84120 207600 84150
rect 207900 84350 208000 84380
rect 207900 84150 207910 84350
rect 207980 84150 208000 84350
rect 207900 84120 208000 84150
rect 196000 84100 196120 84120
rect 196380 84100 196620 84120
rect 196880 84100 197120 84120
rect 197380 84100 197620 84120
rect 197880 84100 198120 84120
rect 198380 84100 198620 84120
rect 198880 84100 199120 84120
rect 199380 84100 199620 84120
rect 199880 84100 200120 84120
rect 200380 84100 200620 84120
rect 200880 84100 201120 84120
rect 201380 84100 201620 84120
rect 201880 84100 202120 84120
rect 202380 84100 202620 84120
rect 202880 84100 203120 84120
rect 203380 84100 203620 84120
rect 203880 84100 204120 84120
rect 204380 84100 204620 84120
rect 204880 84100 205120 84120
rect 205380 84100 205620 84120
rect 205880 84100 206120 84120
rect 206380 84100 206620 84120
rect 206880 84100 207120 84120
rect 207380 84100 207620 84120
rect 207880 84100 208000 84120
rect 196000 84090 208000 84100
rect 196000 84020 196150 84090
rect 196350 84020 196650 84090
rect 196850 84020 197150 84090
rect 197350 84020 197650 84090
rect 197850 84020 198150 84090
rect 198350 84020 198650 84090
rect 198850 84020 199150 84090
rect 199350 84020 199650 84090
rect 199850 84020 200150 84090
rect 200350 84020 200650 84090
rect 200850 84020 201150 84090
rect 201350 84020 201650 84090
rect 201850 84020 202150 84090
rect 202350 84020 202650 84090
rect 202850 84020 203150 84090
rect 203350 84020 203650 84090
rect 203850 84020 204150 84090
rect 204350 84020 204650 84090
rect 204850 84020 205150 84090
rect 205350 84020 205650 84090
rect 205850 84020 206150 84090
rect 206350 84020 206650 84090
rect 206850 84020 207150 84090
rect 207350 84020 207650 84090
rect 207850 84020 208000 84090
rect 196000 83980 208000 84020
rect 196000 83910 196150 83980
rect 196350 83910 196650 83980
rect 196850 83910 197150 83980
rect 197350 83910 197650 83980
rect 197850 83910 198150 83980
rect 198350 83910 198650 83980
rect 198850 83910 199150 83980
rect 199350 83910 199650 83980
rect 199850 83910 200150 83980
rect 200350 83910 200650 83980
rect 200850 83910 201150 83980
rect 201350 83910 201650 83980
rect 201850 83910 202150 83980
rect 202350 83910 202650 83980
rect 202850 83910 203150 83980
rect 203350 83910 203650 83980
rect 203850 83910 204150 83980
rect 204350 83910 204650 83980
rect 204850 83910 205150 83980
rect 205350 83910 205650 83980
rect 205850 83910 206150 83980
rect 206350 83910 206650 83980
rect 206850 83910 207150 83980
rect 207350 83910 207650 83980
rect 207850 83910 208000 83980
rect 196000 83900 208000 83910
rect 196000 83880 196120 83900
rect 196380 83880 196620 83900
rect 196880 83880 197120 83900
rect 197380 83880 197620 83900
rect 197880 83880 198120 83900
rect 198380 83880 198620 83900
rect 198880 83880 199120 83900
rect 199380 83880 199620 83900
rect 199880 83880 200120 83900
rect 200380 83880 200620 83900
rect 200880 83880 201120 83900
rect 201380 83880 201620 83900
rect 201880 83880 202120 83900
rect 202380 83880 202620 83900
rect 202880 83880 203120 83900
rect 203380 83880 203620 83900
rect 203880 83880 204120 83900
rect 204380 83880 204620 83900
rect 204880 83880 205120 83900
rect 205380 83880 205620 83900
rect 205880 83880 206120 83900
rect 206380 83880 206620 83900
rect 206880 83880 207120 83900
rect 207380 83880 207620 83900
rect 207880 83880 208000 83900
rect 196000 83850 196100 83880
rect 196000 83650 196020 83850
rect 196090 83650 196100 83850
rect 196000 83620 196100 83650
rect 196400 83850 196600 83880
rect 196400 83650 196410 83850
rect 196480 83650 196520 83850
rect 196590 83650 196600 83850
rect 196400 83620 196600 83650
rect 196900 83850 197100 83880
rect 196900 83650 196910 83850
rect 196980 83650 197020 83850
rect 197090 83650 197100 83850
rect 196900 83620 197100 83650
rect 197400 83850 197600 83880
rect 197400 83650 197410 83850
rect 197480 83650 197520 83850
rect 197590 83650 197600 83850
rect 197400 83620 197600 83650
rect 197900 83850 198100 83880
rect 197900 83650 197910 83850
rect 197980 83650 198020 83850
rect 198090 83650 198100 83850
rect 197900 83620 198100 83650
rect 198400 83850 198600 83880
rect 198400 83650 198410 83850
rect 198480 83650 198520 83850
rect 198590 83650 198600 83850
rect 198400 83620 198600 83650
rect 198900 83850 199100 83880
rect 198900 83650 198910 83850
rect 198980 83650 199020 83850
rect 199090 83650 199100 83850
rect 198900 83620 199100 83650
rect 199400 83850 199600 83880
rect 199400 83650 199410 83850
rect 199480 83650 199520 83850
rect 199590 83650 199600 83850
rect 199400 83620 199600 83650
rect 199900 83850 200100 83880
rect 199900 83650 199910 83850
rect 199980 83650 200020 83850
rect 200090 83650 200100 83850
rect 199900 83620 200100 83650
rect 200400 83850 200600 83880
rect 200400 83650 200410 83850
rect 200480 83650 200520 83850
rect 200590 83650 200600 83850
rect 200400 83620 200600 83650
rect 200900 83850 201100 83880
rect 200900 83650 200910 83850
rect 200980 83650 201020 83850
rect 201090 83650 201100 83850
rect 200900 83620 201100 83650
rect 201400 83850 201600 83880
rect 201400 83650 201410 83850
rect 201480 83650 201520 83850
rect 201590 83650 201600 83850
rect 201400 83620 201600 83650
rect 201900 83850 202100 83880
rect 201900 83650 201910 83850
rect 201980 83650 202020 83850
rect 202090 83650 202100 83850
rect 201900 83620 202100 83650
rect 202400 83850 202600 83880
rect 202400 83650 202410 83850
rect 202480 83650 202520 83850
rect 202590 83650 202600 83850
rect 202400 83620 202600 83650
rect 202900 83850 203100 83880
rect 202900 83650 202910 83850
rect 202980 83650 203020 83850
rect 203090 83650 203100 83850
rect 202900 83620 203100 83650
rect 203400 83850 203600 83880
rect 203400 83650 203410 83850
rect 203480 83650 203520 83850
rect 203590 83650 203600 83850
rect 203400 83620 203600 83650
rect 203900 83850 204100 83880
rect 203900 83650 203910 83850
rect 203980 83650 204020 83850
rect 204090 83650 204100 83850
rect 203900 83620 204100 83650
rect 204400 83850 204600 83880
rect 204400 83650 204410 83850
rect 204480 83650 204520 83850
rect 204590 83650 204600 83850
rect 204400 83620 204600 83650
rect 204900 83850 205100 83880
rect 204900 83650 204910 83850
rect 204980 83650 205020 83850
rect 205090 83650 205100 83850
rect 204900 83620 205100 83650
rect 205400 83850 205600 83880
rect 205400 83650 205410 83850
rect 205480 83650 205520 83850
rect 205590 83650 205600 83850
rect 205400 83620 205600 83650
rect 205900 83850 206100 83880
rect 205900 83650 205910 83850
rect 205980 83650 206020 83850
rect 206090 83650 206100 83850
rect 205900 83620 206100 83650
rect 206400 83850 206600 83880
rect 206400 83650 206410 83850
rect 206480 83650 206520 83850
rect 206590 83650 206600 83850
rect 206400 83620 206600 83650
rect 206900 83850 207100 83880
rect 206900 83650 206910 83850
rect 206980 83650 207020 83850
rect 207090 83650 207100 83850
rect 206900 83620 207100 83650
rect 207400 83850 207600 83880
rect 207400 83650 207410 83850
rect 207480 83650 207520 83850
rect 207590 83650 207600 83850
rect 207400 83620 207600 83650
rect 207900 83850 208000 83880
rect 207900 83650 207910 83850
rect 207980 83650 208000 83850
rect 207900 83620 208000 83650
rect 196000 83600 196120 83620
rect 196380 83600 196620 83620
rect 196880 83600 197120 83620
rect 197380 83600 197620 83620
rect 197880 83600 198120 83620
rect 198380 83600 198620 83620
rect 198880 83600 199120 83620
rect 199380 83600 199620 83620
rect 199880 83600 200120 83620
rect 200380 83600 200620 83620
rect 200880 83600 201120 83620
rect 201380 83600 201620 83620
rect 201880 83600 202120 83620
rect 202380 83600 202620 83620
rect 202880 83600 203120 83620
rect 203380 83600 203620 83620
rect 203880 83600 204120 83620
rect 204380 83600 204620 83620
rect 204880 83600 205120 83620
rect 205380 83600 205620 83620
rect 205880 83600 206120 83620
rect 206380 83600 206620 83620
rect 206880 83600 207120 83620
rect 207380 83600 207620 83620
rect 207880 83600 208000 83620
rect 196000 83590 208000 83600
rect 196000 83520 196150 83590
rect 196350 83520 196650 83590
rect 196850 83520 197150 83590
rect 197350 83520 197650 83590
rect 197850 83520 198150 83590
rect 198350 83520 198650 83590
rect 198850 83520 199150 83590
rect 199350 83520 199650 83590
rect 199850 83520 200150 83590
rect 200350 83520 200650 83590
rect 200850 83520 201150 83590
rect 201350 83520 201650 83590
rect 201850 83520 202150 83590
rect 202350 83520 202650 83590
rect 202850 83520 203150 83590
rect 203350 83520 203650 83590
rect 203850 83520 204150 83590
rect 204350 83520 204650 83590
rect 204850 83520 205150 83590
rect 205350 83520 205650 83590
rect 205850 83520 206150 83590
rect 206350 83520 206650 83590
rect 206850 83520 207150 83590
rect 207350 83520 207650 83590
rect 207850 83520 208000 83590
rect 196000 83480 208000 83520
rect 196000 83410 196150 83480
rect 196350 83410 196650 83480
rect 196850 83410 197150 83480
rect 197350 83410 197650 83480
rect 197850 83410 198150 83480
rect 198350 83410 198650 83480
rect 198850 83410 199150 83480
rect 199350 83410 199650 83480
rect 199850 83410 200150 83480
rect 200350 83410 200650 83480
rect 200850 83410 201150 83480
rect 201350 83410 201650 83480
rect 201850 83410 202150 83480
rect 202350 83410 202650 83480
rect 202850 83410 203150 83480
rect 203350 83410 203650 83480
rect 203850 83410 204150 83480
rect 204350 83410 204650 83480
rect 204850 83410 205150 83480
rect 205350 83410 205650 83480
rect 205850 83410 206150 83480
rect 206350 83410 206650 83480
rect 206850 83410 207150 83480
rect 207350 83410 207650 83480
rect 207850 83410 208000 83480
rect 196000 83400 208000 83410
rect 196000 83380 196120 83400
rect 196380 83380 196620 83400
rect 196880 83380 197120 83400
rect 197380 83380 197620 83400
rect 197880 83380 198120 83400
rect 198380 83380 198620 83400
rect 198880 83380 199120 83400
rect 199380 83380 199620 83400
rect 199880 83380 200120 83400
rect 200380 83380 200620 83400
rect 200880 83380 201120 83400
rect 201380 83380 201620 83400
rect 201880 83380 202120 83400
rect 202380 83380 202620 83400
rect 202880 83380 203120 83400
rect 203380 83380 203620 83400
rect 203880 83380 204120 83400
rect 204380 83380 204620 83400
rect 204880 83380 205120 83400
rect 205380 83380 205620 83400
rect 205880 83380 206120 83400
rect 206380 83380 206620 83400
rect 206880 83380 207120 83400
rect 207380 83380 207620 83400
rect 207880 83380 208000 83400
rect 196000 83350 196100 83380
rect 196000 83150 196020 83350
rect 196090 83150 196100 83350
rect 196000 83120 196100 83150
rect 196400 83350 196600 83380
rect 196400 83150 196410 83350
rect 196480 83150 196520 83350
rect 196590 83150 196600 83350
rect 196400 83120 196600 83150
rect 196900 83350 197100 83380
rect 196900 83150 196910 83350
rect 196980 83150 197020 83350
rect 197090 83150 197100 83350
rect 196900 83120 197100 83150
rect 197400 83350 197600 83380
rect 197400 83150 197410 83350
rect 197480 83150 197520 83350
rect 197590 83150 197600 83350
rect 197400 83120 197600 83150
rect 197900 83350 198100 83380
rect 197900 83150 197910 83350
rect 197980 83150 198020 83350
rect 198090 83150 198100 83350
rect 197900 83120 198100 83150
rect 198400 83350 198600 83380
rect 198400 83150 198410 83350
rect 198480 83150 198520 83350
rect 198590 83150 198600 83350
rect 198400 83120 198600 83150
rect 198900 83350 199100 83380
rect 198900 83150 198910 83350
rect 198980 83150 199020 83350
rect 199090 83150 199100 83350
rect 198900 83120 199100 83150
rect 199400 83350 199600 83380
rect 199400 83150 199410 83350
rect 199480 83150 199520 83350
rect 199590 83150 199600 83350
rect 199400 83120 199600 83150
rect 199900 83350 200100 83380
rect 199900 83150 199910 83350
rect 199980 83150 200020 83350
rect 200090 83150 200100 83350
rect 199900 83120 200100 83150
rect 200400 83350 200600 83380
rect 200400 83150 200410 83350
rect 200480 83150 200520 83350
rect 200590 83150 200600 83350
rect 200400 83120 200600 83150
rect 200900 83350 201100 83380
rect 200900 83150 200910 83350
rect 200980 83150 201020 83350
rect 201090 83150 201100 83350
rect 200900 83120 201100 83150
rect 201400 83350 201600 83380
rect 201400 83150 201410 83350
rect 201480 83150 201520 83350
rect 201590 83150 201600 83350
rect 201400 83120 201600 83150
rect 201900 83350 202100 83380
rect 201900 83150 201910 83350
rect 201980 83150 202020 83350
rect 202090 83150 202100 83350
rect 201900 83120 202100 83150
rect 202400 83350 202600 83380
rect 202400 83150 202410 83350
rect 202480 83150 202520 83350
rect 202590 83150 202600 83350
rect 202400 83120 202600 83150
rect 202900 83350 203100 83380
rect 202900 83150 202910 83350
rect 202980 83150 203020 83350
rect 203090 83150 203100 83350
rect 202900 83120 203100 83150
rect 203400 83350 203600 83380
rect 203400 83150 203410 83350
rect 203480 83150 203520 83350
rect 203590 83150 203600 83350
rect 203400 83120 203600 83150
rect 203900 83350 204100 83380
rect 203900 83150 203910 83350
rect 203980 83150 204020 83350
rect 204090 83150 204100 83350
rect 203900 83120 204100 83150
rect 204400 83350 204600 83380
rect 204400 83150 204410 83350
rect 204480 83150 204520 83350
rect 204590 83150 204600 83350
rect 204400 83120 204600 83150
rect 204900 83350 205100 83380
rect 204900 83150 204910 83350
rect 204980 83150 205020 83350
rect 205090 83150 205100 83350
rect 204900 83120 205100 83150
rect 205400 83350 205600 83380
rect 205400 83150 205410 83350
rect 205480 83150 205520 83350
rect 205590 83150 205600 83350
rect 205400 83120 205600 83150
rect 205900 83350 206100 83380
rect 205900 83150 205910 83350
rect 205980 83150 206020 83350
rect 206090 83150 206100 83350
rect 205900 83120 206100 83150
rect 206400 83350 206600 83380
rect 206400 83150 206410 83350
rect 206480 83150 206520 83350
rect 206590 83150 206600 83350
rect 206400 83120 206600 83150
rect 206900 83350 207100 83380
rect 206900 83150 206910 83350
rect 206980 83150 207020 83350
rect 207090 83150 207100 83350
rect 206900 83120 207100 83150
rect 207400 83350 207600 83380
rect 207400 83150 207410 83350
rect 207480 83150 207520 83350
rect 207590 83150 207600 83350
rect 207400 83120 207600 83150
rect 207900 83350 208000 83380
rect 207900 83150 207910 83350
rect 207980 83150 208000 83350
rect 207900 83120 208000 83150
rect 196000 83100 196120 83120
rect 196380 83100 196620 83120
rect 196880 83100 197120 83120
rect 197380 83100 197620 83120
rect 197880 83100 198120 83120
rect 198380 83100 198620 83120
rect 198880 83100 199120 83120
rect 199380 83100 199620 83120
rect 199880 83100 200120 83120
rect 200380 83100 200620 83120
rect 200880 83100 201120 83120
rect 201380 83100 201620 83120
rect 201880 83100 202120 83120
rect 202380 83100 202620 83120
rect 202880 83100 203120 83120
rect 203380 83100 203620 83120
rect 203880 83100 204120 83120
rect 204380 83100 204620 83120
rect 204880 83100 205120 83120
rect 205380 83100 205620 83120
rect 205880 83100 206120 83120
rect 206380 83100 206620 83120
rect 206880 83100 207120 83120
rect 207380 83100 207620 83120
rect 207880 83100 208000 83120
rect 196000 83090 208000 83100
rect 196000 83020 196150 83090
rect 196350 83020 196650 83090
rect 196850 83020 197150 83090
rect 197350 83020 197650 83090
rect 197850 83020 198150 83090
rect 198350 83020 198650 83090
rect 198850 83020 199150 83090
rect 199350 83020 199650 83090
rect 199850 83020 200150 83090
rect 200350 83020 200650 83090
rect 200850 83020 201150 83090
rect 201350 83020 201650 83090
rect 201850 83020 202150 83090
rect 202350 83020 202650 83090
rect 202850 83020 203150 83090
rect 203350 83020 203650 83090
rect 203850 83020 204150 83090
rect 204350 83020 204650 83090
rect 204850 83020 205150 83090
rect 205350 83020 205650 83090
rect 205850 83020 206150 83090
rect 206350 83020 206650 83090
rect 206850 83020 207150 83090
rect 207350 83020 207650 83090
rect 207850 83020 208000 83090
rect 196000 82980 208000 83020
rect 196000 82910 196150 82980
rect 196350 82910 196650 82980
rect 196850 82910 197150 82980
rect 197350 82910 197650 82980
rect 197850 82910 198150 82980
rect 198350 82910 198650 82980
rect 198850 82910 199150 82980
rect 199350 82910 199650 82980
rect 199850 82910 200150 82980
rect 200350 82910 200650 82980
rect 200850 82910 201150 82980
rect 201350 82910 201650 82980
rect 201850 82910 202150 82980
rect 202350 82910 202650 82980
rect 202850 82910 203150 82980
rect 203350 82910 203650 82980
rect 203850 82910 204150 82980
rect 204350 82910 204650 82980
rect 204850 82910 205150 82980
rect 205350 82910 205650 82980
rect 205850 82910 206150 82980
rect 206350 82910 206650 82980
rect 206850 82910 207150 82980
rect 207350 82910 207650 82980
rect 207850 82910 208000 82980
rect 196000 82900 208000 82910
rect 196000 82880 196120 82900
rect 196380 82880 196620 82900
rect 196880 82880 197120 82900
rect 197380 82880 197620 82900
rect 197880 82880 198120 82900
rect 198380 82880 198620 82900
rect 198880 82880 199120 82900
rect 199380 82880 199620 82900
rect 199880 82880 200120 82900
rect 200380 82880 200620 82900
rect 200880 82880 201120 82900
rect 201380 82880 201620 82900
rect 201880 82880 202120 82900
rect 202380 82880 202620 82900
rect 202880 82880 203120 82900
rect 203380 82880 203620 82900
rect 203880 82880 204120 82900
rect 204380 82880 204620 82900
rect 204880 82880 205120 82900
rect 205380 82880 205620 82900
rect 205880 82880 206120 82900
rect 206380 82880 206620 82900
rect 206880 82880 207120 82900
rect 207380 82880 207620 82900
rect 207880 82880 208000 82900
rect 196000 82850 196100 82880
rect 196000 82650 196020 82850
rect 196090 82650 196100 82850
rect 196000 82620 196100 82650
rect 196400 82850 196600 82880
rect 196400 82650 196410 82850
rect 196480 82650 196520 82850
rect 196590 82650 196600 82850
rect 196400 82620 196600 82650
rect 196900 82850 197100 82880
rect 196900 82650 196910 82850
rect 196980 82650 197020 82850
rect 197090 82650 197100 82850
rect 196900 82620 197100 82650
rect 197400 82850 197600 82880
rect 197400 82650 197410 82850
rect 197480 82650 197520 82850
rect 197590 82650 197600 82850
rect 197400 82620 197600 82650
rect 197900 82850 198100 82880
rect 197900 82650 197910 82850
rect 197980 82650 198020 82850
rect 198090 82650 198100 82850
rect 197900 82620 198100 82650
rect 198400 82850 198600 82880
rect 198400 82650 198410 82850
rect 198480 82650 198520 82850
rect 198590 82650 198600 82850
rect 198400 82620 198600 82650
rect 198900 82850 199100 82880
rect 198900 82650 198910 82850
rect 198980 82650 199020 82850
rect 199090 82650 199100 82850
rect 198900 82620 199100 82650
rect 199400 82850 199600 82880
rect 199400 82650 199410 82850
rect 199480 82650 199520 82850
rect 199590 82650 199600 82850
rect 199400 82620 199600 82650
rect 199900 82850 200100 82880
rect 199900 82650 199910 82850
rect 199980 82650 200020 82850
rect 200090 82650 200100 82850
rect 199900 82620 200100 82650
rect 200400 82850 200600 82880
rect 200400 82650 200410 82850
rect 200480 82650 200520 82850
rect 200590 82650 200600 82850
rect 200400 82620 200600 82650
rect 200900 82850 201100 82880
rect 200900 82650 200910 82850
rect 200980 82650 201020 82850
rect 201090 82650 201100 82850
rect 200900 82620 201100 82650
rect 201400 82850 201600 82880
rect 201400 82650 201410 82850
rect 201480 82650 201520 82850
rect 201590 82650 201600 82850
rect 201400 82620 201600 82650
rect 201900 82850 202100 82880
rect 201900 82650 201910 82850
rect 201980 82650 202020 82850
rect 202090 82650 202100 82850
rect 201900 82620 202100 82650
rect 202400 82850 202600 82880
rect 202400 82650 202410 82850
rect 202480 82650 202520 82850
rect 202590 82650 202600 82850
rect 202400 82620 202600 82650
rect 202900 82850 203100 82880
rect 202900 82650 202910 82850
rect 202980 82650 203020 82850
rect 203090 82650 203100 82850
rect 202900 82620 203100 82650
rect 203400 82850 203600 82880
rect 203400 82650 203410 82850
rect 203480 82650 203520 82850
rect 203590 82650 203600 82850
rect 203400 82620 203600 82650
rect 203900 82850 204100 82880
rect 203900 82650 203910 82850
rect 203980 82650 204020 82850
rect 204090 82650 204100 82850
rect 203900 82620 204100 82650
rect 204400 82850 204600 82880
rect 204400 82650 204410 82850
rect 204480 82650 204520 82850
rect 204590 82650 204600 82850
rect 204400 82620 204600 82650
rect 204900 82850 205100 82880
rect 204900 82650 204910 82850
rect 204980 82650 205020 82850
rect 205090 82650 205100 82850
rect 204900 82620 205100 82650
rect 205400 82850 205600 82880
rect 205400 82650 205410 82850
rect 205480 82650 205520 82850
rect 205590 82650 205600 82850
rect 205400 82620 205600 82650
rect 205900 82850 206100 82880
rect 205900 82650 205910 82850
rect 205980 82650 206020 82850
rect 206090 82650 206100 82850
rect 205900 82620 206100 82650
rect 206400 82850 206600 82880
rect 206400 82650 206410 82850
rect 206480 82650 206520 82850
rect 206590 82650 206600 82850
rect 206400 82620 206600 82650
rect 206900 82850 207100 82880
rect 206900 82650 206910 82850
rect 206980 82650 207020 82850
rect 207090 82650 207100 82850
rect 206900 82620 207100 82650
rect 207400 82850 207600 82880
rect 207400 82650 207410 82850
rect 207480 82650 207520 82850
rect 207590 82650 207600 82850
rect 207400 82620 207600 82650
rect 207900 82850 208000 82880
rect 207900 82650 207910 82850
rect 207980 82650 208000 82850
rect 207900 82620 208000 82650
rect 196000 82600 196120 82620
rect 196380 82600 196620 82620
rect 196880 82600 197120 82620
rect 197380 82600 197620 82620
rect 197880 82600 198120 82620
rect 198380 82600 198620 82620
rect 198880 82600 199120 82620
rect 199380 82600 199620 82620
rect 199880 82600 200120 82620
rect 200380 82600 200620 82620
rect 200880 82600 201120 82620
rect 201380 82600 201620 82620
rect 201880 82600 202120 82620
rect 202380 82600 202620 82620
rect 202880 82600 203120 82620
rect 203380 82600 203620 82620
rect 203880 82600 204120 82620
rect 204380 82600 204620 82620
rect 204880 82600 205120 82620
rect 205380 82600 205620 82620
rect 205880 82600 206120 82620
rect 206380 82600 206620 82620
rect 206880 82600 207120 82620
rect 207380 82600 207620 82620
rect 207880 82600 208000 82620
rect 196000 82590 208000 82600
rect 196000 82520 196150 82590
rect 196350 82520 196650 82590
rect 196850 82520 197150 82590
rect 197350 82520 197650 82590
rect 197850 82520 198150 82590
rect 198350 82520 198650 82590
rect 198850 82520 199150 82590
rect 199350 82520 199650 82590
rect 199850 82520 200150 82590
rect 200350 82520 200650 82590
rect 200850 82520 201150 82590
rect 201350 82520 201650 82590
rect 201850 82520 202150 82590
rect 202350 82520 202650 82590
rect 202850 82520 203150 82590
rect 203350 82520 203650 82590
rect 203850 82520 204150 82590
rect 204350 82520 204650 82590
rect 204850 82520 205150 82590
rect 205350 82520 205650 82590
rect 205850 82520 206150 82590
rect 206350 82520 206650 82590
rect 206850 82520 207150 82590
rect 207350 82520 207650 82590
rect 207850 82520 208000 82590
rect 196000 82480 208000 82520
rect 196000 82410 196150 82480
rect 196350 82410 196650 82480
rect 196850 82410 197150 82480
rect 197350 82410 197650 82480
rect 197850 82410 198150 82480
rect 198350 82410 198650 82480
rect 198850 82410 199150 82480
rect 199350 82410 199650 82480
rect 199850 82410 200150 82480
rect 200350 82410 200650 82480
rect 200850 82410 201150 82480
rect 201350 82410 201650 82480
rect 201850 82410 202150 82480
rect 202350 82410 202650 82480
rect 202850 82410 203150 82480
rect 203350 82410 203650 82480
rect 203850 82410 204150 82480
rect 204350 82410 204650 82480
rect 204850 82410 205150 82480
rect 205350 82410 205650 82480
rect 205850 82410 206150 82480
rect 206350 82410 206650 82480
rect 206850 82410 207150 82480
rect 207350 82410 207650 82480
rect 207850 82410 208000 82480
rect 196000 82400 208000 82410
rect 196000 82380 196120 82400
rect 196380 82380 196620 82400
rect 196880 82380 197120 82400
rect 197380 82380 197620 82400
rect 197880 82380 198120 82400
rect 198380 82380 198620 82400
rect 198880 82380 199120 82400
rect 199380 82380 199620 82400
rect 199880 82380 200120 82400
rect 200380 82380 200620 82400
rect 200880 82380 201120 82400
rect 201380 82380 201620 82400
rect 201880 82380 202120 82400
rect 202380 82380 202620 82400
rect 202880 82380 203120 82400
rect 203380 82380 203620 82400
rect 203880 82380 204120 82400
rect 204380 82380 204620 82400
rect 204880 82380 205120 82400
rect 205380 82380 205620 82400
rect 205880 82380 206120 82400
rect 206380 82380 206620 82400
rect 206880 82380 207120 82400
rect 207380 82380 207620 82400
rect 207880 82380 208000 82400
rect 196000 82350 196100 82380
rect 196000 82150 196020 82350
rect 196090 82150 196100 82350
rect 196000 82120 196100 82150
rect 196400 82350 196600 82380
rect 196400 82150 196410 82350
rect 196480 82150 196520 82350
rect 196590 82150 196600 82350
rect 196400 82120 196600 82150
rect 196900 82350 197100 82380
rect 196900 82150 196910 82350
rect 196980 82150 197020 82350
rect 197090 82150 197100 82350
rect 196900 82120 197100 82150
rect 197400 82350 197600 82380
rect 197400 82150 197410 82350
rect 197480 82150 197520 82350
rect 197590 82150 197600 82350
rect 197400 82120 197600 82150
rect 197900 82350 198100 82380
rect 197900 82150 197910 82350
rect 197980 82150 198020 82350
rect 198090 82150 198100 82350
rect 197900 82120 198100 82150
rect 198400 82350 198600 82380
rect 198400 82150 198410 82350
rect 198480 82150 198520 82350
rect 198590 82150 198600 82350
rect 198400 82120 198600 82150
rect 198900 82350 199100 82380
rect 198900 82150 198910 82350
rect 198980 82150 199020 82350
rect 199090 82150 199100 82350
rect 198900 82120 199100 82150
rect 199400 82350 199600 82380
rect 199400 82150 199410 82350
rect 199480 82150 199520 82350
rect 199590 82150 199600 82350
rect 199400 82120 199600 82150
rect 199900 82350 200100 82380
rect 199900 82150 199910 82350
rect 199980 82150 200020 82350
rect 200090 82150 200100 82350
rect 199900 82120 200100 82150
rect 200400 82350 200600 82380
rect 200400 82150 200410 82350
rect 200480 82150 200520 82350
rect 200590 82150 200600 82350
rect 200400 82120 200600 82150
rect 200900 82350 201100 82380
rect 200900 82150 200910 82350
rect 200980 82150 201020 82350
rect 201090 82150 201100 82350
rect 200900 82120 201100 82150
rect 201400 82350 201600 82380
rect 201400 82150 201410 82350
rect 201480 82150 201520 82350
rect 201590 82150 201600 82350
rect 201400 82120 201600 82150
rect 201900 82350 202100 82380
rect 201900 82150 201910 82350
rect 201980 82150 202020 82350
rect 202090 82150 202100 82350
rect 201900 82120 202100 82150
rect 202400 82350 202600 82380
rect 202400 82150 202410 82350
rect 202480 82150 202520 82350
rect 202590 82150 202600 82350
rect 202400 82120 202600 82150
rect 202900 82350 203100 82380
rect 202900 82150 202910 82350
rect 202980 82150 203020 82350
rect 203090 82150 203100 82350
rect 202900 82120 203100 82150
rect 203400 82350 203600 82380
rect 203400 82150 203410 82350
rect 203480 82150 203520 82350
rect 203590 82150 203600 82350
rect 203400 82120 203600 82150
rect 203900 82350 204100 82380
rect 203900 82150 203910 82350
rect 203980 82150 204020 82350
rect 204090 82150 204100 82350
rect 203900 82120 204100 82150
rect 204400 82350 204600 82380
rect 204400 82150 204410 82350
rect 204480 82150 204520 82350
rect 204590 82150 204600 82350
rect 204400 82120 204600 82150
rect 204900 82350 205100 82380
rect 204900 82150 204910 82350
rect 204980 82150 205020 82350
rect 205090 82150 205100 82350
rect 204900 82120 205100 82150
rect 205400 82350 205600 82380
rect 205400 82150 205410 82350
rect 205480 82150 205520 82350
rect 205590 82150 205600 82350
rect 205400 82120 205600 82150
rect 205900 82350 206100 82380
rect 205900 82150 205910 82350
rect 205980 82150 206020 82350
rect 206090 82150 206100 82350
rect 205900 82120 206100 82150
rect 206400 82350 206600 82380
rect 206400 82150 206410 82350
rect 206480 82150 206520 82350
rect 206590 82150 206600 82350
rect 206400 82120 206600 82150
rect 206900 82350 207100 82380
rect 206900 82150 206910 82350
rect 206980 82150 207020 82350
rect 207090 82150 207100 82350
rect 206900 82120 207100 82150
rect 207400 82350 207600 82380
rect 207400 82150 207410 82350
rect 207480 82150 207520 82350
rect 207590 82150 207600 82350
rect 207400 82120 207600 82150
rect 207900 82350 208000 82380
rect 207900 82150 207910 82350
rect 207980 82150 208000 82350
rect 207900 82120 208000 82150
rect 196000 82100 196120 82120
rect 196380 82100 196620 82120
rect 196880 82100 197120 82120
rect 197380 82100 197620 82120
rect 197880 82100 198120 82120
rect 198380 82100 198620 82120
rect 198880 82100 199120 82120
rect 199380 82100 199620 82120
rect 199880 82100 200120 82120
rect 200380 82100 200620 82120
rect 200880 82100 201120 82120
rect 201380 82100 201620 82120
rect 201880 82100 202120 82120
rect 202380 82100 202620 82120
rect 202880 82100 203120 82120
rect 203380 82100 203620 82120
rect 203880 82100 204120 82120
rect 204380 82100 204620 82120
rect 204880 82100 205120 82120
rect 205380 82100 205620 82120
rect 205880 82100 206120 82120
rect 206380 82100 206620 82120
rect 206880 82100 207120 82120
rect 207380 82100 207620 82120
rect 207880 82100 208000 82120
rect 196000 82090 208000 82100
rect 196000 82020 196150 82090
rect 196350 82020 196650 82090
rect 196850 82020 197150 82090
rect 197350 82020 197650 82090
rect 197850 82020 198150 82090
rect 198350 82020 198650 82090
rect 198850 82020 199150 82090
rect 199350 82020 199650 82090
rect 199850 82020 200150 82090
rect 200350 82020 200650 82090
rect 200850 82020 201150 82090
rect 201350 82020 201650 82090
rect 201850 82020 202150 82090
rect 202350 82020 202650 82090
rect 202850 82020 203150 82090
rect 203350 82020 203650 82090
rect 203850 82020 204150 82090
rect 204350 82020 204650 82090
rect 204850 82020 205150 82090
rect 205350 82020 205650 82090
rect 205850 82020 206150 82090
rect 206350 82020 206650 82090
rect 206850 82020 207150 82090
rect 207350 82020 207650 82090
rect 207850 82020 208000 82090
rect 196000 81980 208000 82020
rect 196000 81910 196150 81980
rect 196350 81910 196650 81980
rect 196850 81910 197150 81980
rect 197350 81910 197650 81980
rect 197850 81910 198150 81980
rect 198350 81910 198650 81980
rect 198850 81910 199150 81980
rect 199350 81910 199650 81980
rect 199850 81910 200150 81980
rect 200350 81910 200650 81980
rect 200850 81910 201150 81980
rect 201350 81910 201650 81980
rect 201850 81910 202150 81980
rect 202350 81910 202650 81980
rect 202850 81910 203150 81980
rect 203350 81910 203650 81980
rect 203850 81910 204150 81980
rect 204350 81910 204650 81980
rect 204850 81910 205150 81980
rect 205350 81910 205650 81980
rect 205850 81910 206150 81980
rect 206350 81910 206650 81980
rect 206850 81910 207150 81980
rect 207350 81910 207650 81980
rect 207850 81910 208000 81980
rect 196000 81900 208000 81910
rect 196000 81880 196120 81900
rect 196380 81880 196620 81900
rect 196880 81880 197120 81900
rect 197380 81880 197620 81900
rect 197880 81880 198120 81900
rect 198380 81880 198620 81900
rect 198880 81880 199120 81900
rect 199380 81880 199620 81900
rect 199880 81880 200120 81900
rect 200380 81880 200620 81900
rect 200880 81880 201120 81900
rect 201380 81880 201620 81900
rect 201880 81880 202120 81900
rect 202380 81880 202620 81900
rect 202880 81880 203120 81900
rect 203380 81880 203620 81900
rect 203880 81880 204120 81900
rect 204380 81880 204620 81900
rect 204880 81880 205120 81900
rect 205380 81880 205620 81900
rect 205880 81880 206120 81900
rect 206380 81880 206620 81900
rect 206880 81880 207120 81900
rect 207380 81880 207620 81900
rect 207880 81880 208000 81900
rect 196000 81850 196100 81880
rect 196000 81650 196020 81850
rect 196090 81650 196100 81850
rect 196000 81620 196100 81650
rect 196400 81850 196600 81880
rect 196400 81650 196410 81850
rect 196480 81650 196520 81850
rect 196590 81650 196600 81850
rect 196400 81620 196600 81650
rect 196900 81850 197100 81880
rect 196900 81650 196910 81850
rect 196980 81650 197020 81850
rect 197090 81650 197100 81850
rect 196900 81620 197100 81650
rect 197400 81850 197600 81880
rect 197400 81650 197410 81850
rect 197480 81650 197520 81850
rect 197590 81650 197600 81850
rect 197400 81620 197600 81650
rect 197900 81850 198100 81880
rect 197900 81650 197910 81850
rect 197980 81650 198020 81850
rect 198090 81650 198100 81850
rect 197900 81620 198100 81650
rect 198400 81850 198600 81880
rect 198400 81650 198410 81850
rect 198480 81650 198520 81850
rect 198590 81650 198600 81850
rect 198400 81620 198600 81650
rect 198900 81850 199100 81880
rect 198900 81650 198910 81850
rect 198980 81650 199020 81850
rect 199090 81650 199100 81850
rect 198900 81620 199100 81650
rect 199400 81850 199600 81880
rect 199400 81650 199410 81850
rect 199480 81650 199520 81850
rect 199590 81650 199600 81850
rect 199400 81620 199600 81650
rect 199900 81850 200100 81880
rect 199900 81650 199910 81850
rect 199980 81650 200020 81850
rect 200090 81650 200100 81850
rect 199900 81620 200100 81650
rect 200400 81850 200600 81880
rect 200400 81650 200410 81850
rect 200480 81650 200520 81850
rect 200590 81650 200600 81850
rect 200400 81620 200600 81650
rect 200900 81850 201100 81880
rect 200900 81650 200910 81850
rect 200980 81650 201020 81850
rect 201090 81650 201100 81850
rect 200900 81620 201100 81650
rect 201400 81850 201600 81880
rect 201400 81650 201410 81850
rect 201480 81650 201520 81850
rect 201590 81650 201600 81850
rect 201400 81620 201600 81650
rect 201900 81850 202100 81880
rect 201900 81650 201910 81850
rect 201980 81650 202020 81850
rect 202090 81650 202100 81850
rect 201900 81620 202100 81650
rect 202400 81850 202600 81880
rect 202400 81650 202410 81850
rect 202480 81650 202520 81850
rect 202590 81650 202600 81850
rect 202400 81620 202600 81650
rect 202900 81850 203100 81880
rect 202900 81650 202910 81850
rect 202980 81650 203020 81850
rect 203090 81650 203100 81850
rect 202900 81620 203100 81650
rect 203400 81850 203600 81880
rect 203400 81650 203410 81850
rect 203480 81650 203520 81850
rect 203590 81650 203600 81850
rect 203400 81620 203600 81650
rect 203900 81850 204100 81880
rect 203900 81650 203910 81850
rect 203980 81650 204020 81850
rect 204090 81650 204100 81850
rect 203900 81620 204100 81650
rect 204400 81850 204600 81880
rect 204400 81650 204410 81850
rect 204480 81650 204520 81850
rect 204590 81650 204600 81850
rect 204400 81620 204600 81650
rect 204900 81850 205100 81880
rect 204900 81650 204910 81850
rect 204980 81650 205020 81850
rect 205090 81650 205100 81850
rect 204900 81620 205100 81650
rect 205400 81850 205600 81880
rect 205400 81650 205410 81850
rect 205480 81650 205520 81850
rect 205590 81650 205600 81850
rect 205400 81620 205600 81650
rect 205900 81850 206100 81880
rect 205900 81650 205910 81850
rect 205980 81650 206020 81850
rect 206090 81650 206100 81850
rect 205900 81620 206100 81650
rect 206400 81850 206600 81880
rect 206400 81650 206410 81850
rect 206480 81650 206520 81850
rect 206590 81650 206600 81850
rect 206400 81620 206600 81650
rect 206900 81850 207100 81880
rect 206900 81650 206910 81850
rect 206980 81650 207020 81850
rect 207090 81650 207100 81850
rect 206900 81620 207100 81650
rect 207400 81850 207600 81880
rect 207400 81650 207410 81850
rect 207480 81650 207520 81850
rect 207590 81650 207600 81850
rect 207400 81620 207600 81650
rect 207900 81850 208000 81880
rect 207900 81650 207910 81850
rect 207980 81650 208000 81850
rect 207900 81620 208000 81650
rect 196000 81600 196120 81620
rect 196380 81600 196620 81620
rect 196880 81600 197120 81620
rect 197380 81600 197620 81620
rect 197880 81600 198120 81620
rect 198380 81600 198620 81620
rect 198880 81600 199120 81620
rect 199380 81600 199620 81620
rect 199880 81600 200120 81620
rect 200380 81600 200620 81620
rect 200880 81600 201120 81620
rect 201380 81600 201620 81620
rect 201880 81600 202120 81620
rect 202380 81600 202620 81620
rect 202880 81600 203120 81620
rect 203380 81600 203620 81620
rect 203880 81600 204120 81620
rect 204380 81600 204620 81620
rect 204880 81600 205120 81620
rect 205380 81600 205620 81620
rect 205880 81600 206120 81620
rect 206380 81600 206620 81620
rect 206880 81600 207120 81620
rect 207380 81600 207620 81620
rect 207880 81600 208000 81620
rect 196000 81590 208000 81600
rect 196000 81520 196150 81590
rect 196350 81520 196650 81590
rect 196850 81520 197150 81590
rect 197350 81520 197650 81590
rect 197850 81520 198150 81590
rect 198350 81520 198650 81590
rect 198850 81520 199150 81590
rect 199350 81520 199650 81590
rect 199850 81520 200150 81590
rect 200350 81520 200650 81590
rect 200850 81520 201150 81590
rect 201350 81520 201650 81590
rect 201850 81520 202150 81590
rect 202350 81520 202650 81590
rect 202850 81520 203150 81590
rect 203350 81520 203650 81590
rect 203850 81520 204150 81590
rect 204350 81520 204650 81590
rect 204850 81520 205150 81590
rect 205350 81520 205650 81590
rect 205850 81520 206150 81590
rect 206350 81520 206650 81590
rect 206850 81520 207150 81590
rect 207350 81520 207650 81590
rect 207850 81520 208000 81590
rect 196000 81480 208000 81520
rect 196000 81410 196150 81480
rect 196350 81410 196650 81480
rect 196850 81410 197150 81480
rect 197350 81410 197650 81480
rect 197850 81410 198150 81480
rect 198350 81410 198650 81480
rect 198850 81410 199150 81480
rect 199350 81410 199650 81480
rect 199850 81410 200150 81480
rect 200350 81410 200650 81480
rect 200850 81410 201150 81480
rect 201350 81410 201650 81480
rect 201850 81410 202150 81480
rect 202350 81410 202650 81480
rect 202850 81410 203150 81480
rect 203350 81410 203650 81480
rect 203850 81410 204150 81480
rect 204350 81410 204650 81480
rect 204850 81410 205150 81480
rect 205350 81410 205650 81480
rect 205850 81410 206150 81480
rect 206350 81410 206650 81480
rect 206850 81410 207150 81480
rect 207350 81410 207650 81480
rect 207850 81410 208000 81480
rect 196000 81400 208000 81410
rect 196000 81380 196120 81400
rect 196380 81380 196620 81400
rect 196880 81380 197120 81400
rect 197380 81380 197620 81400
rect 197880 81380 198120 81400
rect 198380 81380 198620 81400
rect 198880 81380 199120 81400
rect 199380 81380 199620 81400
rect 199880 81380 200120 81400
rect 200380 81380 200620 81400
rect 200880 81380 201120 81400
rect 201380 81380 201620 81400
rect 201880 81380 202120 81400
rect 202380 81380 202620 81400
rect 202880 81380 203120 81400
rect 203380 81380 203620 81400
rect 203880 81380 204120 81400
rect 204380 81380 204620 81400
rect 204880 81380 205120 81400
rect 205380 81380 205620 81400
rect 205880 81380 206120 81400
rect 206380 81380 206620 81400
rect 206880 81380 207120 81400
rect 207380 81380 207620 81400
rect 207880 81380 208000 81400
rect 196000 81350 196100 81380
rect 196000 81150 196020 81350
rect 196090 81150 196100 81350
rect 196000 81120 196100 81150
rect 196400 81350 196600 81380
rect 196400 81150 196410 81350
rect 196480 81150 196520 81350
rect 196590 81150 196600 81350
rect 196400 81120 196600 81150
rect 196900 81350 197100 81380
rect 196900 81150 196910 81350
rect 196980 81150 197020 81350
rect 197090 81150 197100 81350
rect 196900 81120 197100 81150
rect 197400 81350 197600 81380
rect 197400 81150 197410 81350
rect 197480 81150 197520 81350
rect 197590 81150 197600 81350
rect 197400 81120 197600 81150
rect 197900 81350 198100 81380
rect 197900 81150 197910 81350
rect 197980 81150 198020 81350
rect 198090 81150 198100 81350
rect 197900 81120 198100 81150
rect 198400 81350 198600 81380
rect 198400 81150 198410 81350
rect 198480 81150 198520 81350
rect 198590 81150 198600 81350
rect 198400 81120 198600 81150
rect 198900 81350 199100 81380
rect 198900 81150 198910 81350
rect 198980 81150 199020 81350
rect 199090 81150 199100 81350
rect 198900 81120 199100 81150
rect 199400 81350 199600 81380
rect 199400 81150 199410 81350
rect 199480 81150 199520 81350
rect 199590 81150 199600 81350
rect 199400 81120 199600 81150
rect 199900 81350 200100 81380
rect 199900 81150 199910 81350
rect 199980 81150 200020 81350
rect 200090 81150 200100 81350
rect 199900 81120 200100 81150
rect 200400 81350 200600 81380
rect 200400 81150 200410 81350
rect 200480 81150 200520 81350
rect 200590 81150 200600 81350
rect 200400 81120 200600 81150
rect 200900 81350 201100 81380
rect 200900 81150 200910 81350
rect 200980 81150 201020 81350
rect 201090 81150 201100 81350
rect 200900 81120 201100 81150
rect 201400 81350 201600 81380
rect 201400 81150 201410 81350
rect 201480 81150 201520 81350
rect 201590 81150 201600 81350
rect 201400 81120 201600 81150
rect 201900 81350 202100 81380
rect 201900 81150 201910 81350
rect 201980 81150 202020 81350
rect 202090 81150 202100 81350
rect 201900 81120 202100 81150
rect 202400 81350 202600 81380
rect 202400 81150 202410 81350
rect 202480 81150 202520 81350
rect 202590 81150 202600 81350
rect 202400 81120 202600 81150
rect 202900 81350 203100 81380
rect 202900 81150 202910 81350
rect 202980 81150 203020 81350
rect 203090 81150 203100 81350
rect 202900 81120 203100 81150
rect 203400 81350 203600 81380
rect 203400 81150 203410 81350
rect 203480 81150 203520 81350
rect 203590 81150 203600 81350
rect 203400 81120 203600 81150
rect 203900 81350 204100 81380
rect 203900 81150 203910 81350
rect 203980 81150 204020 81350
rect 204090 81150 204100 81350
rect 203900 81120 204100 81150
rect 204400 81350 204600 81380
rect 204400 81150 204410 81350
rect 204480 81150 204520 81350
rect 204590 81150 204600 81350
rect 204400 81120 204600 81150
rect 204900 81350 205100 81380
rect 204900 81150 204910 81350
rect 204980 81150 205020 81350
rect 205090 81150 205100 81350
rect 204900 81120 205100 81150
rect 205400 81350 205600 81380
rect 205400 81150 205410 81350
rect 205480 81150 205520 81350
rect 205590 81150 205600 81350
rect 205400 81120 205600 81150
rect 205900 81350 206100 81380
rect 205900 81150 205910 81350
rect 205980 81150 206020 81350
rect 206090 81150 206100 81350
rect 205900 81120 206100 81150
rect 206400 81350 206600 81380
rect 206400 81150 206410 81350
rect 206480 81150 206520 81350
rect 206590 81150 206600 81350
rect 206400 81120 206600 81150
rect 206900 81350 207100 81380
rect 206900 81150 206910 81350
rect 206980 81150 207020 81350
rect 207090 81150 207100 81350
rect 206900 81120 207100 81150
rect 207400 81350 207600 81380
rect 207400 81150 207410 81350
rect 207480 81150 207520 81350
rect 207590 81150 207600 81350
rect 207400 81120 207600 81150
rect 207900 81350 208000 81380
rect 207900 81150 207910 81350
rect 207980 81150 208000 81350
rect 207900 81120 208000 81150
rect 196000 81100 196120 81120
rect 196380 81100 196620 81120
rect 196880 81100 197120 81120
rect 197380 81100 197620 81120
rect 197880 81100 198120 81120
rect 198380 81100 198620 81120
rect 198880 81100 199120 81120
rect 199380 81100 199620 81120
rect 199880 81100 200120 81120
rect 200380 81100 200620 81120
rect 200880 81100 201120 81120
rect 201380 81100 201620 81120
rect 201880 81100 202120 81120
rect 202380 81100 202620 81120
rect 202880 81100 203120 81120
rect 203380 81100 203620 81120
rect 203880 81100 204120 81120
rect 204380 81100 204620 81120
rect 204880 81100 205120 81120
rect 205380 81100 205620 81120
rect 205880 81100 206120 81120
rect 206380 81100 206620 81120
rect 206880 81100 207120 81120
rect 207380 81100 207620 81120
rect 207880 81100 208000 81120
rect 196000 81090 208000 81100
rect 196000 81020 196150 81090
rect 196350 81020 196650 81090
rect 196850 81020 197150 81090
rect 197350 81020 197650 81090
rect 197850 81020 198150 81090
rect 198350 81020 198650 81090
rect 198850 81020 199150 81090
rect 199350 81020 199650 81090
rect 199850 81020 200150 81090
rect 200350 81020 200650 81090
rect 200850 81020 201150 81090
rect 201350 81020 201650 81090
rect 201850 81020 202150 81090
rect 202350 81020 202650 81090
rect 202850 81020 203150 81090
rect 203350 81020 203650 81090
rect 203850 81020 204150 81090
rect 204350 81020 204650 81090
rect 204850 81020 205150 81090
rect 205350 81020 205650 81090
rect 205850 81020 206150 81090
rect 206350 81020 206650 81090
rect 206850 81020 207150 81090
rect 207350 81020 207650 81090
rect 207850 81020 208000 81090
rect 196000 80980 208000 81020
rect 196000 80910 196150 80980
rect 196350 80910 196650 80980
rect 196850 80910 197150 80980
rect 197350 80910 197650 80980
rect 197850 80910 198150 80980
rect 198350 80910 198650 80980
rect 198850 80910 199150 80980
rect 199350 80910 199650 80980
rect 199850 80910 200150 80980
rect 200350 80910 200650 80980
rect 200850 80910 201150 80980
rect 201350 80910 201650 80980
rect 201850 80910 202150 80980
rect 202350 80910 202650 80980
rect 202850 80910 203150 80980
rect 203350 80910 203650 80980
rect 203850 80910 204150 80980
rect 204350 80910 204650 80980
rect 204850 80910 205150 80980
rect 205350 80910 205650 80980
rect 205850 80910 206150 80980
rect 206350 80910 206650 80980
rect 206850 80910 207150 80980
rect 207350 80910 207650 80980
rect 207850 80910 208000 80980
rect 196000 80900 208000 80910
rect 196000 80880 196120 80900
rect 196380 80880 196620 80900
rect 196880 80880 197120 80900
rect 197380 80880 197620 80900
rect 197880 80880 198120 80900
rect 198380 80880 198620 80900
rect 198880 80880 199120 80900
rect 199380 80880 199620 80900
rect 199880 80880 200120 80900
rect 200380 80880 200620 80900
rect 200880 80880 201120 80900
rect 201380 80880 201620 80900
rect 201880 80880 202120 80900
rect 202380 80880 202620 80900
rect 202880 80880 203120 80900
rect 203380 80880 203620 80900
rect 203880 80880 204120 80900
rect 204380 80880 204620 80900
rect 204880 80880 205120 80900
rect 205380 80880 205620 80900
rect 205880 80880 206120 80900
rect 206380 80880 206620 80900
rect 206880 80880 207120 80900
rect 207380 80880 207620 80900
rect 207880 80880 208000 80900
rect 196000 80850 196100 80880
rect 196000 80650 196020 80850
rect 196090 80650 196100 80850
rect 196000 80620 196100 80650
rect 196400 80850 196600 80880
rect 196400 80650 196410 80850
rect 196480 80650 196520 80850
rect 196590 80650 196600 80850
rect 196400 80620 196600 80650
rect 196900 80850 197100 80880
rect 196900 80650 196910 80850
rect 196980 80650 197020 80850
rect 197090 80650 197100 80850
rect 196900 80620 197100 80650
rect 197400 80850 197600 80880
rect 197400 80650 197410 80850
rect 197480 80650 197520 80850
rect 197590 80650 197600 80850
rect 197400 80620 197600 80650
rect 197900 80850 198100 80880
rect 197900 80650 197910 80850
rect 197980 80650 198020 80850
rect 198090 80650 198100 80850
rect 197900 80620 198100 80650
rect 198400 80850 198600 80880
rect 198400 80650 198410 80850
rect 198480 80650 198520 80850
rect 198590 80650 198600 80850
rect 198400 80620 198600 80650
rect 198900 80850 199100 80880
rect 198900 80650 198910 80850
rect 198980 80650 199020 80850
rect 199090 80650 199100 80850
rect 198900 80620 199100 80650
rect 199400 80850 199600 80880
rect 199400 80650 199410 80850
rect 199480 80650 199520 80850
rect 199590 80650 199600 80850
rect 199400 80620 199600 80650
rect 199900 80850 200100 80880
rect 199900 80650 199910 80850
rect 199980 80650 200020 80850
rect 200090 80650 200100 80850
rect 199900 80620 200100 80650
rect 200400 80850 200600 80880
rect 200400 80650 200410 80850
rect 200480 80650 200520 80850
rect 200590 80650 200600 80850
rect 200400 80620 200600 80650
rect 200900 80850 201100 80880
rect 200900 80650 200910 80850
rect 200980 80650 201020 80850
rect 201090 80650 201100 80850
rect 200900 80620 201100 80650
rect 201400 80850 201600 80880
rect 201400 80650 201410 80850
rect 201480 80650 201520 80850
rect 201590 80650 201600 80850
rect 201400 80620 201600 80650
rect 201900 80850 202100 80880
rect 201900 80650 201910 80850
rect 201980 80650 202020 80850
rect 202090 80650 202100 80850
rect 201900 80620 202100 80650
rect 202400 80850 202600 80880
rect 202400 80650 202410 80850
rect 202480 80650 202520 80850
rect 202590 80650 202600 80850
rect 202400 80620 202600 80650
rect 202900 80850 203100 80880
rect 202900 80650 202910 80850
rect 202980 80650 203020 80850
rect 203090 80650 203100 80850
rect 202900 80620 203100 80650
rect 203400 80850 203600 80880
rect 203400 80650 203410 80850
rect 203480 80650 203520 80850
rect 203590 80650 203600 80850
rect 203400 80620 203600 80650
rect 203900 80850 204100 80880
rect 203900 80650 203910 80850
rect 203980 80650 204020 80850
rect 204090 80650 204100 80850
rect 203900 80620 204100 80650
rect 204400 80850 204600 80880
rect 204400 80650 204410 80850
rect 204480 80650 204520 80850
rect 204590 80650 204600 80850
rect 204400 80620 204600 80650
rect 204900 80850 205100 80880
rect 204900 80650 204910 80850
rect 204980 80650 205020 80850
rect 205090 80650 205100 80850
rect 204900 80620 205100 80650
rect 205400 80850 205600 80880
rect 205400 80650 205410 80850
rect 205480 80650 205520 80850
rect 205590 80650 205600 80850
rect 205400 80620 205600 80650
rect 205900 80850 206100 80880
rect 205900 80650 205910 80850
rect 205980 80650 206020 80850
rect 206090 80650 206100 80850
rect 205900 80620 206100 80650
rect 206400 80850 206600 80880
rect 206400 80650 206410 80850
rect 206480 80650 206520 80850
rect 206590 80650 206600 80850
rect 206400 80620 206600 80650
rect 206900 80850 207100 80880
rect 206900 80650 206910 80850
rect 206980 80650 207020 80850
rect 207090 80650 207100 80850
rect 206900 80620 207100 80650
rect 207400 80850 207600 80880
rect 207400 80650 207410 80850
rect 207480 80650 207520 80850
rect 207590 80650 207600 80850
rect 207400 80620 207600 80650
rect 207900 80850 208000 80880
rect 207900 80650 207910 80850
rect 207980 80650 208000 80850
rect 207900 80620 208000 80650
rect 196000 80600 196120 80620
rect 196380 80600 196620 80620
rect 196880 80600 197120 80620
rect 197380 80600 197620 80620
rect 197880 80600 198120 80620
rect 198380 80600 198620 80620
rect 198880 80600 199120 80620
rect 199380 80600 199620 80620
rect 199880 80600 200120 80620
rect 200380 80600 200620 80620
rect 200880 80600 201120 80620
rect 201380 80600 201620 80620
rect 201880 80600 202120 80620
rect 202380 80600 202620 80620
rect 202880 80600 203120 80620
rect 203380 80600 203620 80620
rect 203880 80600 204120 80620
rect 204380 80600 204620 80620
rect 204880 80600 205120 80620
rect 205380 80600 205620 80620
rect 205880 80600 206120 80620
rect 206380 80600 206620 80620
rect 206880 80600 207120 80620
rect 207380 80600 207620 80620
rect 207880 80600 208000 80620
rect 196000 80590 208000 80600
rect 196000 80520 196150 80590
rect 196350 80520 196650 80590
rect 196850 80520 197150 80590
rect 197350 80520 197650 80590
rect 197850 80520 198150 80590
rect 198350 80520 198650 80590
rect 198850 80520 199150 80590
rect 199350 80520 199650 80590
rect 199850 80520 200150 80590
rect 200350 80520 200650 80590
rect 200850 80520 201150 80590
rect 201350 80520 201650 80590
rect 201850 80520 202150 80590
rect 202350 80520 202650 80590
rect 202850 80520 203150 80590
rect 203350 80520 203650 80590
rect 203850 80520 204150 80590
rect 204350 80520 204650 80590
rect 204850 80520 205150 80590
rect 205350 80520 205650 80590
rect 205850 80520 206150 80590
rect 206350 80520 206650 80590
rect 206850 80520 207150 80590
rect 207350 80520 207650 80590
rect 207850 80520 208000 80590
rect 196000 80480 208000 80520
rect 196000 80410 196150 80480
rect 196350 80410 196650 80480
rect 196850 80410 197150 80480
rect 197350 80410 197650 80480
rect 197850 80410 198150 80480
rect 198350 80410 198650 80480
rect 198850 80410 199150 80480
rect 199350 80410 199650 80480
rect 199850 80410 200150 80480
rect 200350 80410 200650 80480
rect 200850 80410 201150 80480
rect 201350 80410 201650 80480
rect 201850 80410 202150 80480
rect 202350 80410 202650 80480
rect 202850 80410 203150 80480
rect 203350 80410 203650 80480
rect 203850 80410 204150 80480
rect 204350 80410 204650 80480
rect 204850 80410 205150 80480
rect 205350 80410 205650 80480
rect 205850 80410 206150 80480
rect 206350 80410 206650 80480
rect 206850 80410 207150 80480
rect 207350 80410 207650 80480
rect 207850 80410 208000 80480
rect 196000 80400 208000 80410
rect 196000 80380 196120 80400
rect 196380 80380 196620 80400
rect 196880 80380 197120 80400
rect 197380 80380 197620 80400
rect 197880 80380 198120 80400
rect 198380 80380 198620 80400
rect 198880 80380 199120 80400
rect 199380 80380 199620 80400
rect 199880 80380 200120 80400
rect 200380 80380 200620 80400
rect 200880 80380 201120 80400
rect 201380 80380 201620 80400
rect 201880 80380 202120 80400
rect 202380 80380 202620 80400
rect 202880 80380 203120 80400
rect 203380 80380 203620 80400
rect 203880 80380 204120 80400
rect 204380 80380 204620 80400
rect 204880 80380 205120 80400
rect 205380 80380 205620 80400
rect 205880 80380 206120 80400
rect 206380 80380 206620 80400
rect 206880 80380 207120 80400
rect 207380 80380 207620 80400
rect 207880 80380 208000 80400
rect 196000 80350 196100 80380
rect 196000 80150 196020 80350
rect 196090 80150 196100 80350
rect 196000 80120 196100 80150
rect 196400 80350 196600 80380
rect 196400 80150 196410 80350
rect 196480 80150 196520 80350
rect 196590 80150 196600 80350
rect 196400 80120 196600 80150
rect 196900 80350 197100 80380
rect 196900 80150 196910 80350
rect 196980 80150 197020 80350
rect 197090 80150 197100 80350
rect 196900 80120 197100 80150
rect 197400 80350 197600 80380
rect 197400 80150 197410 80350
rect 197480 80150 197520 80350
rect 197590 80150 197600 80350
rect 197400 80120 197600 80150
rect 197900 80350 198100 80380
rect 197900 80150 197910 80350
rect 197980 80150 198020 80350
rect 198090 80150 198100 80350
rect 197900 80120 198100 80150
rect 198400 80350 198600 80380
rect 198400 80150 198410 80350
rect 198480 80150 198520 80350
rect 198590 80150 198600 80350
rect 198400 80120 198600 80150
rect 198900 80350 199100 80380
rect 198900 80150 198910 80350
rect 198980 80150 199020 80350
rect 199090 80150 199100 80350
rect 198900 80120 199100 80150
rect 199400 80350 199600 80380
rect 199400 80150 199410 80350
rect 199480 80150 199520 80350
rect 199590 80150 199600 80350
rect 199400 80120 199600 80150
rect 199900 80350 200100 80380
rect 199900 80150 199910 80350
rect 199980 80150 200020 80350
rect 200090 80150 200100 80350
rect 199900 80120 200100 80150
rect 200400 80350 200600 80380
rect 200400 80150 200410 80350
rect 200480 80150 200520 80350
rect 200590 80150 200600 80350
rect 200400 80120 200600 80150
rect 200900 80350 201100 80380
rect 200900 80150 200910 80350
rect 200980 80150 201020 80350
rect 201090 80150 201100 80350
rect 200900 80120 201100 80150
rect 201400 80350 201600 80380
rect 201400 80150 201410 80350
rect 201480 80150 201520 80350
rect 201590 80150 201600 80350
rect 201400 80120 201600 80150
rect 201900 80350 202100 80380
rect 201900 80150 201910 80350
rect 201980 80150 202020 80350
rect 202090 80150 202100 80350
rect 201900 80120 202100 80150
rect 202400 80350 202600 80380
rect 202400 80150 202410 80350
rect 202480 80150 202520 80350
rect 202590 80150 202600 80350
rect 202400 80120 202600 80150
rect 202900 80350 203100 80380
rect 202900 80150 202910 80350
rect 202980 80150 203020 80350
rect 203090 80150 203100 80350
rect 202900 80120 203100 80150
rect 203400 80350 203600 80380
rect 203400 80150 203410 80350
rect 203480 80150 203520 80350
rect 203590 80150 203600 80350
rect 203400 80120 203600 80150
rect 203900 80350 204100 80380
rect 203900 80150 203910 80350
rect 203980 80150 204020 80350
rect 204090 80150 204100 80350
rect 203900 80120 204100 80150
rect 204400 80350 204600 80380
rect 204400 80150 204410 80350
rect 204480 80150 204520 80350
rect 204590 80150 204600 80350
rect 204400 80120 204600 80150
rect 204900 80350 205100 80380
rect 204900 80150 204910 80350
rect 204980 80150 205020 80350
rect 205090 80150 205100 80350
rect 204900 80120 205100 80150
rect 205400 80350 205600 80380
rect 205400 80150 205410 80350
rect 205480 80150 205520 80350
rect 205590 80150 205600 80350
rect 205400 80120 205600 80150
rect 205900 80350 206100 80380
rect 205900 80150 205910 80350
rect 205980 80150 206020 80350
rect 206090 80150 206100 80350
rect 205900 80120 206100 80150
rect 206400 80350 206600 80380
rect 206400 80150 206410 80350
rect 206480 80150 206520 80350
rect 206590 80150 206600 80350
rect 206400 80120 206600 80150
rect 206900 80350 207100 80380
rect 206900 80150 206910 80350
rect 206980 80150 207020 80350
rect 207090 80150 207100 80350
rect 206900 80120 207100 80150
rect 207400 80350 207600 80380
rect 207400 80150 207410 80350
rect 207480 80150 207520 80350
rect 207590 80150 207600 80350
rect 207400 80120 207600 80150
rect 207900 80350 208000 80380
rect 207900 80150 207910 80350
rect 207980 80150 208000 80350
rect 207900 80120 208000 80150
rect 196000 80100 196120 80120
rect 196380 80100 196620 80120
rect 196880 80100 197120 80120
rect 197380 80100 197620 80120
rect 197880 80100 198120 80120
rect 198380 80100 198620 80120
rect 198880 80100 199120 80120
rect 199380 80100 199620 80120
rect 199880 80100 200120 80120
rect 200380 80100 200620 80120
rect 200880 80100 201120 80120
rect 201380 80100 201620 80120
rect 201880 80100 202120 80120
rect 202380 80100 202620 80120
rect 202880 80100 203120 80120
rect 203380 80100 203620 80120
rect 203880 80100 204120 80120
rect 204380 80100 204620 80120
rect 204880 80100 205120 80120
rect 205380 80100 205620 80120
rect 205880 80100 206120 80120
rect 206380 80100 206620 80120
rect 206880 80100 207120 80120
rect 207380 80100 207620 80120
rect 207880 80100 208000 80120
rect 196000 80090 208000 80100
rect 196000 80020 196150 80090
rect 196350 80020 196650 80090
rect 196850 80020 197150 80090
rect 197350 80020 197650 80090
rect 197850 80020 198150 80090
rect 198350 80020 198650 80090
rect 198850 80020 199150 80090
rect 199350 80020 199650 80090
rect 199850 80020 200150 80090
rect 200350 80020 200650 80090
rect 200850 80020 201150 80090
rect 201350 80020 201650 80090
rect 201850 80020 202150 80090
rect 202350 80020 202650 80090
rect 202850 80020 203150 80090
rect 203350 80020 203650 80090
rect 203850 80020 204150 80090
rect 204350 80020 204650 80090
rect 204850 80020 205150 80090
rect 205350 80020 205650 80090
rect 205850 80020 206150 80090
rect 206350 80020 206650 80090
rect 206850 80020 207150 80090
rect 207350 80020 207650 80090
rect 207850 80020 208000 80090
rect 196000 79980 208000 80020
rect 196000 79910 196150 79980
rect 196350 79910 196650 79980
rect 196850 79910 197150 79980
rect 197350 79910 197650 79980
rect 197850 79910 198150 79980
rect 198350 79910 198650 79980
rect 198850 79910 199150 79980
rect 199350 79910 199650 79980
rect 199850 79910 200150 79980
rect 200350 79910 200650 79980
rect 200850 79910 201150 79980
rect 201350 79910 201650 79980
rect 201850 79910 202150 79980
rect 202350 79910 202650 79980
rect 202850 79910 203150 79980
rect 203350 79910 203650 79980
rect 203850 79910 204150 79980
rect 204350 79910 204650 79980
rect 204850 79910 205150 79980
rect 205350 79910 205650 79980
rect 205850 79910 206150 79980
rect 206350 79910 206650 79980
rect 206850 79910 207150 79980
rect 207350 79910 207650 79980
rect 207850 79910 208000 79980
rect 196000 79900 208000 79910
rect 196000 79880 196120 79900
rect 196380 79880 196620 79900
rect 196880 79880 197120 79900
rect 197380 79880 197620 79900
rect 197880 79880 198120 79900
rect 198380 79880 198620 79900
rect 198880 79880 199120 79900
rect 199380 79880 199620 79900
rect 199880 79880 200120 79900
rect 200380 79880 200620 79900
rect 200880 79880 201120 79900
rect 201380 79880 201620 79900
rect 201880 79880 202120 79900
rect 202380 79880 202620 79900
rect 202880 79880 203120 79900
rect 203380 79880 203620 79900
rect 203880 79880 204120 79900
rect 204380 79880 204620 79900
rect 204880 79880 205120 79900
rect 205380 79880 205620 79900
rect 205880 79880 206120 79900
rect 206380 79880 206620 79900
rect 206880 79880 207120 79900
rect 207380 79880 207620 79900
rect 207880 79880 208000 79900
rect 196000 79850 196100 79880
rect 196000 79650 196020 79850
rect 196090 79650 196100 79850
rect 196000 79620 196100 79650
rect 196400 79850 196600 79880
rect 196400 79650 196410 79850
rect 196480 79650 196520 79850
rect 196590 79650 196600 79850
rect 196400 79620 196600 79650
rect 196900 79850 197100 79880
rect 196900 79650 196910 79850
rect 196980 79650 197020 79850
rect 197090 79650 197100 79850
rect 196900 79620 197100 79650
rect 197400 79850 197600 79880
rect 197400 79650 197410 79850
rect 197480 79650 197520 79850
rect 197590 79650 197600 79850
rect 197400 79620 197600 79650
rect 197900 79850 198100 79880
rect 197900 79650 197910 79850
rect 197980 79650 198020 79850
rect 198090 79650 198100 79850
rect 197900 79620 198100 79650
rect 198400 79850 198600 79880
rect 198400 79650 198410 79850
rect 198480 79650 198520 79850
rect 198590 79650 198600 79850
rect 198400 79620 198600 79650
rect 198900 79850 199100 79880
rect 198900 79650 198910 79850
rect 198980 79650 199020 79850
rect 199090 79650 199100 79850
rect 198900 79620 199100 79650
rect 199400 79850 199600 79880
rect 199400 79650 199410 79850
rect 199480 79650 199520 79850
rect 199590 79650 199600 79850
rect 199400 79620 199600 79650
rect 199900 79850 200100 79880
rect 199900 79650 199910 79850
rect 199980 79650 200020 79850
rect 200090 79650 200100 79850
rect 199900 79620 200100 79650
rect 200400 79850 200600 79880
rect 200400 79650 200410 79850
rect 200480 79650 200520 79850
rect 200590 79650 200600 79850
rect 200400 79620 200600 79650
rect 200900 79850 201100 79880
rect 200900 79650 200910 79850
rect 200980 79650 201020 79850
rect 201090 79650 201100 79850
rect 200900 79620 201100 79650
rect 201400 79850 201600 79880
rect 201400 79650 201410 79850
rect 201480 79650 201520 79850
rect 201590 79650 201600 79850
rect 201400 79620 201600 79650
rect 201900 79850 202100 79880
rect 201900 79650 201910 79850
rect 201980 79650 202020 79850
rect 202090 79650 202100 79850
rect 201900 79620 202100 79650
rect 202400 79850 202600 79880
rect 202400 79650 202410 79850
rect 202480 79650 202520 79850
rect 202590 79650 202600 79850
rect 202400 79620 202600 79650
rect 202900 79850 203100 79880
rect 202900 79650 202910 79850
rect 202980 79650 203020 79850
rect 203090 79650 203100 79850
rect 202900 79620 203100 79650
rect 203400 79850 203600 79880
rect 203400 79650 203410 79850
rect 203480 79650 203520 79850
rect 203590 79650 203600 79850
rect 203400 79620 203600 79650
rect 203900 79850 204100 79880
rect 203900 79650 203910 79850
rect 203980 79650 204020 79850
rect 204090 79650 204100 79850
rect 203900 79620 204100 79650
rect 204400 79850 204600 79880
rect 204400 79650 204410 79850
rect 204480 79650 204520 79850
rect 204590 79650 204600 79850
rect 204400 79620 204600 79650
rect 204900 79850 205100 79880
rect 204900 79650 204910 79850
rect 204980 79650 205020 79850
rect 205090 79650 205100 79850
rect 204900 79620 205100 79650
rect 205400 79850 205600 79880
rect 205400 79650 205410 79850
rect 205480 79650 205520 79850
rect 205590 79650 205600 79850
rect 205400 79620 205600 79650
rect 205900 79850 206100 79880
rect 205900 79650 205910 79850
rect 205980 79650 206020 79850
rect 206090 79650 206100 79850
rect 205900 79620 206100 79650
rect 206400 79850 206600 79880
rect 206400 79650 206410 79850
rect 206480 79650 206520 79850
rect 206590 79650 206600 79850
rect 206400 79620 206600 79650
rect 206900 79850 207100 79880
rect 206900 79650 206910 79850
rect 206980 79650 207020 79850
rect 207090 79650 207100 79850
rect 206900 79620 207100 79650
rect 207400 79850 207600 79880
rect 207400 79650 207410 79850
rect 207480 79650 207520 79850
rect 207590 79650 207600 79850
rect 207400 79620 207600 79650
rect 207900 79850 208000 79880
rect 207900 79650 207910 79850
rect 207980 79650 208000 79850
rect 207900 79620 208000 79650
rect 196000 79600 196120 79620
rect 196380 79600 196620 79620
rect 196880 79600 197120 79620
rect 197380 79600 197620 79620
rect 197880 79600 198120 79620
rect 198380 79600 198620 79620
rect 198880 79600 199120 79620
rect 199380 79600 199620 79620
rect 199880 79600 200120 79620
rect 200380 79600 200620 79620
rect 200880 79600 201120 79620
rect 201380 79600 201620 79620
rect 201880 79600 202120 79620
rect 202380 79600 202620 79620
rect 202880 79600 203120 79620
rect 203380 79600 203620 79620
rect 203880 79600 204120 79620
rect 204380 79600 204620 79620
rect 204880 79600 205120 79620
rect 205380 79600 205620 79620
rect 205880 79600 206120 79620
rect 206380 79600 206620 79620
rect 206880 79600 207120 79620
rect 207380 79600 207620 79620
rect 207880 79600 208000 79620
rect 196000 79590 208000 79600
rect 196000 79520 196150 79590
rect 196350 79520 196650 79590
rect 196850 79520 197150 79590
rect 197350 79520 197650 79590
rect 197850 79520 198150 79590
rect 198350 79520 198650 79590
rect 198850 79520 199150 79590
rect 199350 79520 199650 79590
rect 199850 79520 200150 79590
rect 200350 79520 200650 79590
rect 200850 79520 201150 79590
rect 201350 79520 201650 79590
rect 201850 79520 202150 79590
rect 202350 79520 202650 79590
rect 202850 79520 203150 79590
rect 203350 79520 203650 79590
rect 203850 79520 204150 79590
rect 204350 79520 204650 79590
rect 204850 79520 205150 79590
rect 205350 79520 205650 79590
rect 205850 79520 206150 79590
rect 206350 79520 206650 79590
rect 206850 79520 207150 79590
rect 207350 79520 207650 79590
rect 207850 79520 208000 79590
rect 196000 79480 208000 79520
rect 196000 79410 196150 79480
rect 196350 79410 196650 79480
rect 196850 79410 197150 79480
rect 197350 79410 197650 79480
rect 197850 79410 198150 79480
rect 198350 79410 198650 79480
rect 198850 79410 199150 79480
rect 199350 79410 199650 79480
rect 199850 79410 200150 79480
rect 200350 79410 200650 79480
rect 200850 79410 201150 79480
rect 201350 79410 201650 79480
rect 201850 79410 202150 79480
rect 202350 79410 202650 79480
rect 202850 79410 203150 79480
rect 203350 79410 203650 79480
rect 203850 79410 204150 79480
rect 204350 79410 204650 79480
rect 204850 79410 205150 79480
rect 205350 79410 205650 79480
rect 205850 79410 206150 79480
rect 206350 79410 206650 79480
rect 206850 79410 207150 79480
rect 207350 79410 207650 79480
rect 207850 79410 208000 79480
rect 196000 79400 208000 79410
rect 196000 79380 196120 79400
rect 196380 79380 196620 79400
rect 196880 79380 197120 79400
rect 197380 79380 197620 79400
rect 197880 79380 198120 79400
rect 198380 79380 198620 79400
rect 198880 79380 199120 79400
rect 199380 79380 199620 79400
rect 199880 79380 200120 79400
rect 200380 79380 200620 79400
rect 200880 79380 201120 79400
rect 201380 79380 201620 79400
rect 201880 79380 202120 79400
rect 202380 79380 202620 79400
rect 202880 79380 203120 79400
rect 203380 79380 203620 79400
rect 203880 79380 204120 79400
rect 204380 79380 204620 79400
rect 204880 79380 205120 79400
rect 205380 79380 205620 79400
rect 205880 79380 206120 79400
rect 206380 79380 206620 79400
rect 206880 79380 207120 79400
rect 207380 79380 207620 79400
rect 207880 79380 208000 79400
rect 196000 79350 196100 79380
rect 196000 79150 196020 79350
rect 196090 79150 196100 79350
rect 196000 79120 196100 79150
rect 196400 79350 196600 79380
rect 196400 79150 196410 79350
rect 196480 79150 196520 79350
rect 196590 79150 196600 79350
rect 196400 79120 196600 79150
rect 196900 79350 197100 79380
rect 196900 79150 196910 79350
rect 196980 79150 197020 79350
rect 197090 79150 197100 79350
rect 196900 79120 197100 79150
rect 197400 79350 197600 79380
rect 197400 79150 197410 79350
rect 197480 79150 197520 79350
rect 197590 79150 197600 79350
rect 197400 79120 197600 79150
rect 197900 79350 198100 79380
rect 197900 79150 197910 79350
rect 197980 79150 198020 79350
rect 198090 79150 198100 79350
rect 197900 79120 198100 79150
rect 198400 79350 198600 79380
rect 198400 79150 198410 79350
rect 198480 79150 198520 79350
rect 198590 79150 198600 79350
rect 198400 79120 198600 79150
rect 198900 79350 199100 79380
rect 198900 79150 198910 79350
rect 198980 79150 199020 79350
rect 199090 79150 199100 79350
rect 198900 79120 199100 79150
rect 199400 79350 199600 79380
rect 199400 79150 199410 79350
rect 199480 79150 199520 79350
rect 199590 79150 199600 79350
rect 199400 79120 199600 79150
rect 199900 79350 200100 79380
rect 199900 79150 199910 79350
rect 199980 79150 200020 79350
rect 200090 79150 200100 79350
rect 199900 79120 200100 79150
rect 200400 79350 200600 79380
rect 200400 79150 200410 79350
rect 200480 79150 200520 79350
rect 200590 79150 200600 79350
rect 200400 79120 200600 79150
rect 200900 79350 201100 79380
rect 200900 79150 200910 79350
rect 200980 79150 201020 79350
rect 201090 79150 201100 79350
rect 200900 79120 201100 79150
rect 201400 79350 201600 79380
rect 201400 79150 201410 79350
rect 201480 79150 201520 79350
rect 201590 79150 201600 79350
rect 201400 79120 201600 79150
rect 201900 79350 202100 79380
rect 201900 79150 201910 79350
rect 201980 79150 202020 79350
rect 202090 79150 202100 79350
rect 201900 79120 202100 79150
rect 202400 79350 202600 79380
rect 202400 79150 202410 79350
rect 202480 79150 202520 79350
rect 202590 79150 202600 79350
rect 202400 79120 202600 79150
rect 202900 79350 203100 79380
rect 202900 79150 202910 79350
rect 202980 79150 203020 79350
rect 203090 79150 203100 79350
rect 202900 79120 203100 79150
rect 203400 79350 203600 79380
rect 203400 79150 203410 79350
rect 203480 79150 203520 79350
rect 203590 79150 203600 79350
rect 203400 79120 203600 79150
rect 203900 79350 204100 79380
rect 203900 79150 203910 79350
rect 203980 79150 204020 79350
rect 204090 79150 204100 79350
rect 203900 79120 204100 79150
rect 204400 79350 204600 79380
rect 204400 79150 204410 79350
rect 204480 79150 204520 79350
rect 204590 79150 204600 79350
rect 204400 79120 204600 79150
rect 204900 79350 205100 79380
rect 204900 79150 204910 79350
rect 204980 79150 205020 79350
rect 205090 79150 205100 79350
rect 204900 79120 205100 79150
rect 205400 79350 205600 79380
rect 205400 79150 205410 79350
rect 205480 79150 205520 79350
rect 205590 79150 205600 79350
rect 205400 79120 205600 79150
rect 205900 79350 206100 79380
rect 205900 79150 205910 79350
rect 205980 79150 206020 79350
rect 206090 79150 206100 79350
rect 205900 79120 206100 79150
rect 206400 79350 206600 79380
rect 206400 79150 206410 79350
rect 206480 79150 206520 79350
rect 206590 79150 206600 79350
rect 206400 79120 206600 79150
rect 206900 79350 207100 79380
rect 206900 79150 206910 79350
rect 206980 79150 207020 79350
rect 207090 79150 207100 79350
rect 206900 79120 207100 79150
rect 207400 79350 207600 79380
rect 207400 79150 207410 79350
rect 207480 79150 207520 79350
rect 207590 79150 207600 79350
rect 207400 79120 207600 79150
rect 207900 79350 208000 79380
rect 207900 79150 207910 79350
rect 207980 79150 208000 79350
rect 207900 79120 208000 79150
rect 196000 79100 196120 79120
rect 196380 79100 196620 79120
rect 196880 79100 197120 79120
rect 197380 79100 197620 79120
rect 197880 79100 198120 79120
rect 198380 79100 198620 79120
rect 198880 79100 199120 79120
rect 199380 79100 199620 79120
rect 199880 79100 200120 79120
rect 200380 79100 200620 79120
rect 200880 79100 201120 79120
rect 201380 79100 201620 79120
rect 201880 79100 202120 79120
rect 202380 79100 202620 79120
rect 202880 79100 203120 79120
rect 203380 79100 203620 79120
rect 203880 79100 204120 79120
rect 204380 79100 204620 79120
rect 204880 79100 205120 79120
rect 205380 79100 205620 79120
rect 205880 79100 206120 79120
rect 206380 79100 206620 79120
rect 206880 79100 207120 79120
rect 207380 79100 207620 79120
rect 207880 79100 208000 79120
rect 196000 79090 208000 79100
rect 196000 79020 196150 79090
rect 196350 79020 196650 79090
rect 196850 79020 197150 79090
rect 197350 79020 197650 79090
rect 197850 79020 198150 79090
rect 198350 79020 198650 79090
rect 198850 79020 199150 79090
rect 199350 79020 199650 79090
rect 199850 79020 200150 79090
rect 200350 79020 200650 79090
rect 200850 79020 201150 79090
rect 201350 79020 201650 79090
rect 201850 79020 202150 79090
rect 202350 79020 202650 79090
rect 202850 79020 203150 79090
rect 203350 79020 203650 79090
rect 203850 79020 204150 79090
rect 204350 79020 204650 79090
rect 204850 79020 205150 79090
rect 205350 79020 205650 79090
rect 205850 79020 206150 79090
rect 206350 79020 206650 79090
rect 206850 79020 207150 79090
rect 207350 79020 207650 79090
rect 207850 79020 208000 79090
rect 196000 78980 208000 79020
rect 196000 78910 196150 78980
rect 196350 78910 196650 78980
rect 196850 78910 197150 78980
rect 197350 78910 197650 78980
rect 197850 78910 198150 78980
rect 198350 78910 198650 78980
rect 198850 78910 199150 78980
rect 199350 78910 199650 78980
rect 199850 78910 200150 78980
rect 200350 78910 200650 78980
rect 200850 78910 201150 78980
rect 201350 78910 201650 78980
rect 201850 78910 202150 78980
rect 202350 78910 202650 78980
rect 202850 78910 203150 78980
rect 203350 78910 203650 78980
rect 203850 78910 204150 78980
rect 204350 78910 204650 78980
rect 204850 78910 205150 78980
rect 205350 78910 205650 78980
rect 205850 78910 206150 78980
rect 206350 78910 206650 78980
rect 206850 78910 207150 78980
rect 207350 78910 207650 78980
rect 207850 78910 208000 78980
rect 196000 78900 208000 78910
rect 196000 78880 196120 78900
rect 196380 78880 196620 78900
rect 196880 78880 197120 78900
rect 197380 78880 197620 78900
rect 197880 78880 198120 78900
rect 198380 78880 198620 78900
rect 198880 78880 199120 78900
rect 199380 78880 199620 78900
rect 199880 78880 200120 78900
rect 200380 78880 200620 78900
rect 200880 78880 201120 78900
rect 201380 78880 201620 78900
rect 201880 78880 202120 78900
rect 202380 78880 202620 78900
rect 202880 78880 203120 78900
rect 203380 78880 203620 78900
rect 203880 78880 204120 78900
rect 204380 78880 204620 78900
rect 204880 78880 205120 78900
rect 205380 78880 205620 78900
rect 205880 78880 206120 78900
rect 206380 78880 206620 78900
rect 206880 78880 207120 78900
rect 207380 78880 207620 78900
rect 207880 78880 208000 78900
rect 196000 78850 196100 78880
rect 196000 78650 196020 78850
rect 196090 78650 196100 78850
rect 196000 78620 196100 78650
rect 196400 78850 196600 78880
rect 196400 78650 196410 78850
rect 196480 78650 196520 78850
rect 196590 78650 196600 78850
rect 196400 78620 196600 78650
rect 196900 78850 197100 78880
rect 196900 78650 196910 78850
rect 196980 78650 197020 78850
rect 197090 78650 197100 78850
rect 196900 78620 197100 78650
rect 197400 78850 197600 78880
rect 197400 78650 197410 78850
rect 197480 78650 197520 78850
rect 197590 78650 197600 78850
rect 197400 78620 197600 78650
rect 197900 78850 198100 78880
rect 197900 78650 197910 78850
rect 197980 78650 198020 78850
rect 198090 78650 198100 78850
rect 197900 78620 198100 78650
rect 198400 78850 198600 78880
rect 198400 78650 198410 78850
rect 198480 78650 198520 78850
rect 198590 78650 198600 78850
rect 198400 78620 198600 78650
rect 198900 78850 199100 78880
rect 198900 78650 198910 78850
rect 198980 78650 199020 78850
rect 199090 78650 199100 78850
rect 198900 78620 199100 78650
rect 199400 78850 199600 78880
rect 199400 78650 199410 78850
rect 199480 78650 199520 78850
rect 199590 78650 199600 78850
rect 199400 78620 199600 78650
rect 199900 78850 200100 78880
rect 199900 78650 199910 78850
rect 199980 78650 200020 78850
rect 200090 78650 200100 78850
rect 199900 78620 200100 78650
rect 200400 78850 200600 78880
rect 200400 78650 200410 78850
rect 200480 78650 200520 78850
rect 200590 78650 200600 78850
rect 200400 78620 200600 78650
rect 200900 78850 201100 78880
rect 200900 78650 200910 78850
rect 200980 78650 201020 78850
rect 201090 78650 201100 78850
rect 200900 78620 201100 78650
rect 201400 78850 201600 78880
rect 201400 78650 201410 78850
rect 201480 78650 201520 78850
rect 201590 78650 201600 78850
rect 201400 78620 201600 78650
rect 201900 78850 202100 78880
rect 201900 78650 201910 78850
rect 201980 78650 202020 78850
rect 202090 78650 202100 78850
rect 201900 78620 202100 78650
rect 202400 78850 202600 78880
rect 202400 78650 202410 78850
rect 202480 78650 202520 78850
rect 202590 78650 202600 78850
rect 202400 78620 202600 78650
rect 202900 78850 203100 78880
rect 202900 78650 202910 78850
rect 202980 78650 203020 78850
rect 203090 78650 203100 78850
rect 202900 78620 203100 78650
rect 203400 78850 203600 78880
rect 203400 78650 203410 78850
rect 203480 78650 203520 78850
rect 203590 78650 203600 78850
rect 203400 78620 203600 78650
rect 203900 78850 204100 78880
rect 203900 78650 203910 78850
rect 203980 78650 204020 78850
rect 204090 78650 204100 78850
rect 203900 78620 204100 78650
rect 204400 78850 204600 78880
rect 204400 78650 204410 78850
rect 204480 78650 204520 78850
rect 204590 78650 204600 78850
rect 204400 78620 204600 78650
rect 204900 78850 205100 78880
rect 204900 78650 204910 78850
rect 204980 78650 205020 78850
rect 205090 78650 205100 78850
rect 204900 78620 205100 78650
rect 205400 78850 205600 78880
rect 205400 78650 205410 78850
rect 205480 78650 205520 78850
rect 205590 78650 205600 78850
rect 205400 78620 205600 78650
rect 205900 78850 206100 78880
rect 205900 78650 205910 78850
rect 205980 78650 206020 78850
rect 206090 78650 206100 78850
rect 205900 78620 206100 78650
rect 206400 78850 206600 78880
rect 206400 78650 206410 78850
rect 206480 78650 206520 78850
rect 206590 78650 206600 78850
rect 206400 78620 206600 78650
rect 206900 78850 207100 78880
rect 206900 78650 206910 78850
rect 206980 78650 207020 78850
rect 207090 78650 207100 78850
rect 206900 78620 207100 78650
rect 207400 78850 207600 78880
rect 207400 78650 207410 78850
rect 207480 78650 207520 78850
rect 207590 78650 207600 78850
rect 207400 78620 207600 78650
rect 207900 78850 208000 78880
rect 207900 78650 207910 78850
rect 207980 78650 208000 78850
rect 207900 78620 208000 78650
rect 196000 78600 196120 78620
rect 196380 78600 196620 78620
rect 196880 78600 197120 78620
rect 197380 78600 197620 78620
rect 197880 78600 198120 78620
rect 198380 78600 198620 78620
rect 198880 78600 199120 78620
rect 199380 78600 199620 78620
rect 199880 78600 200120 78620
rect 200380 78600 200620 78620
rect 200880 78600 201120 78620
rect 201380 78600 201620 78620
rect 201880 78600 202120 78620
rect 202380 78600 202620 78620
rect 202880 78600 203120 78620
rect 203380 78600 203620 78620
rect 203880 78600 204120 78620
rect 204380 78600 204620 78620
rect 204880 78600 205120 78620
rect 205380 78600 205620 78620
rect 205880 78600 206120 78620
rect 206380 78600 206620 78620
rect 206880 78600 207120 78620
rect 207380 78600 207620 78620
rect 207880 78600 208000 78620
rect 196000 78590 208000 78600
rect 196000 78520 196150 78590
rect 196350 78520 196650 78590
rect 196850 78520 197150 78590
rect 197350 78520 197650 78590
rect 197850 78520 198150 78590
rect 198350 78520 198650 78590
rect 198850 78520 199150 78590
rect 199350 78520 199650 78590
rect 199850 78520 200150 78590
rect 200350 78520 200650 78590
rect 200850 78520 201150 78590
rect 201350 78520 201650 78590
rect 201850 78520 202150 78590
rect 202350 78520 202650 78590
rect 202850 78520 203150 78590
rect 203350 78520 203650 78590
rect 203850 78520 204150 78590
rect 204350 78520 204650 78590
rect 204850 78520 205150 78590
rect 205350 78520 205650 78590
rect 205850 78520 206150 78590
rect 206350 78520 206650 78590
rect 206850 78520 207150 78590
rect 207350 78520 207650 78590
rect 207850 78520 208000 78590
rect 196000 78480 208000 78520
rect 196000 78410 196150 78480
rect 196350 78410 196650 78480
rect 196850 78410 197150 78480
rect 197350 78410 197650 78480
rect 197850 78410 198150 78480
rect 198350 78410 198650 78480
rect 198850 78410 199150 78480
rect 199350 78410 199650 78480
rect 199850 78410 200150 78480
rect 200350 78410 200650 78480
rect 200850 78410 201150 78480
rect 201350 78410 201650 78480
rect 201850 78410 202150 78480
rect 202350 78410 202650 78480
rect 202850 78410 203150 78480
rect 203350 78410 203650 78480
rect 203850 78410 204150 78480
rect 204350 78410 204650 78480
rect 204850 78410 205150 78480
rect 205350 78410 205650 78480
rect 205850 78410 206150 78480
rect 206350 78410 206650 78480
rect 206850 78410 207150 78480
rect 207350 78410 207650 78480
rect 207850 78410 208000 78480
rect 196000 78400 208000 78410
rect 196000 78380 196120 78400
rect 196380 78380 196620 78400
rect 196880 78380 197120 78400
rect 197380 78380 197620 78400
rect 197880 78380 198120 78400
rect 198380 78380 198620 78400
rect 198880 78380 199120 78400
rect 199380 78380 199620 78400
rect 199880 78380 200120 78400
rect 200380 78380 200620 78400
rect 200880 78380 201120 78400
rect 201380 78380 201620 78400
rect 201880 78380 202120 78400
rect 202380 78380 202620 78400
rect 202880 78380 203120 78400
rect 203380 78380 203620 78400
rect 203880 78380 204120 78400
rect 204380 78380 204620 78400
rect 204880 78380 205120 78400
rect 205380 78380 205620 78400
rect 205880 78380 206120 78400
rect 206380 78380 206620 78400
rect 206880 78380 207120 78400
rect 207380 78380 207620 78400
rect 207880 78380 208000 78400
rect 196000 78350 196100 78380
rect 196000 78150 196020 78350
rect 196090 78150 196100 78350
rect 196000 78120 196100 78150
rect 196400 78350 196600 78380
rect 196400 78150 196410 78350
rect 196480 78150 196520 78350
rect 196590 78150 196600 78350
rect 196400 78120 196600 78150
rect 196900 78350 197100 78380
rect 196900 78150 196910 78350
rect 196980 78150 197020 78350
rect 197090 78150 197100 78350
rect 196900 78120 197100 78150
rect 197400 78350 197600 78380
rect 197400 78150 197410 78350
rect 197480 78150 197520 78350
rect 197590 78150 197600 78350
rect 197400 78120 197600 78150
rect 197900 78350 198100 78380
rect 197900 78150 197910 78350
rect 197980 78150 198020 78350
rect 198090 78150 198100 78350
rect 197900 78120 198100 78150
rect 198400 78350 198600 78380
rect 198400 78150 198410 78350
rect 198480 78150 198520 78350
rect 198590 78150 198600 78350
rect 198400 78120 198600 78150
rect 198900 78350 199100 78380
rect 198900 78150 198910 78350
rect 198980 78150 199020 78350
rect 199090 78150 199100 78350
rect 198900 78120 199100 78150
rect 199400 78350 199600 78380
rect 199400 78150 199410 78350
rect 199480 78150 199520 78350
rect 199590 78150 199600 78350
rect 199400 78120 199600 78150
rect 199900 78350 200100 78380
rect 199900 78150 199910 78350
rect 199980 78150 200020 78350
rect 200090 78150 200100 78350
rect 199900 78120 200100 78150
rect 200400 78350 200600 78380
rect 200400 78150 200410 78350
rect 200480 78150 200520 78350
rect 200590 78150 200600 78350
rect 200400 78120 200600 78150
rect 200900 78350 201100 78380
rect 200900 78150 200910 78350
rect 200980 78150 201020 78350
rect 201090 78150 201100 78350
rect 200900 78120 201100 78150
rect 201400 78350 201600 78380
rect 201400 78150 201410 78350
rect 201480 78150 201520 78350
rect 201590 78150 201600 78350
rect 201400 78120 201600 78150
rect 201900 78350 202100 78380
rect 201900 78150 201910 78350
rect 201980 78150 202020 78350
rect 202090 78150 202100 78350
rect 201900 78120 202100 78150
rect 202400 78350 202600 78380
rect 202400 78150 202410 78350
rect 202480 78150 202520 78350
rect 202590 78150 202600 78350
rect 202400 78120 202600 78150
rect 202900 78350 203100 78380
rect 202900 78150 202910 78350
rect 202980 78150 203020 78350
rect 203090 78150 203100 78350
rect 202900 78120 203100 78150
rect 203400 78350 203600 78380
rect 203400 78150 203410 78350
rect 203480 78150 203520 78350
rect 203590 78150 203600 78350
rect 203400 78120 203600 78150
rect 203900 78350 204100 78380
rect 203900 78150 203910 78350
rect 203980 78150 204020 78350
rect 204090 78150 204100 78350
rect 203900 78120 204100 78150
rect 204400 78350 204600 78380
rect 204400 78150 204410 78350
rect 204480 78150 204520 78350
rect 204590 78150 204600 78350
rect 204400 78120 204600 78150
rect 204900 78350 205100 78380
rect 204900 78150 204910 78350
rect 204980 78150 205020 78350
rect 205090 78150 205100 78350
rect 204900 78120 205100 78150
rect 205400 78350 205600 78380
rect 205400 78150 205410 78350
rect 205480 78150 205520 78350
rect 205590 78150 205600 78350
rect 205400 78120 205600 78150
rect 205900 78350 206100 78380
rect 205900 78150 205910 78350
rect 205980 78150 206020 78350
rect 206090 78150 206100 78350
rect 205900 78120 206100 78150
rect 206400 78350 206600 78380
rect 206400 78150 206410 78350
rect 206480 78150 206520 78350
rect 206590 78150 206600 78350
rect 206400 78120 206600 78150
rect 206900 78350 207100 78380
rect 206900 78150 206910 78350
rect 206980 78150 207020 78350
rect 207090 78150 207100 78350
rect 206900 78120 207100 78150
rect 207400 78350 207600 78380
rect 207400 78150 207410 78350
rect 207480 78150 207520 78350
rect 207590 78150 207600 78350
rect 207400 78120 207600 78150
rect 207900 78350 208000 78380
rect 207900 78150 207910 78350
rect 207980 78150 208000 78350
rect 207900 78120 208000 78150
rect 196000 78100 196120 78120
rect 196380 78100 196620 78120
rect 196880 78100 197120 78120
rect 197380 78100 197620 78120
rect 197880 78100 198120 78120
rect 198380 78100 198620 78120
rect 198880 78100 199120 78120
rect 199380 78100 199620 78120
rect 199880 78100 200120 78120
rect 200380 78100 200620 78120
rect 200880 78100 201120 78120
rect 201380 78100 201620 78120
rect 201880 78100 202120 78120
rect 202380 78100 202620 78120
rect 202880 78100 203120 78120
rect 203380 78100 203620 78120
rect 203880 78100 204120 78120
rect 204380 78100 204620 78120
rect 204880 78100 205120 78120
rect 205380 78100 205620 78120
rect 205880 78100 206120 78120
rect 206380 78100 206620 78120
rect 206880 78100 207120 78120
rect 207380 78100 207620 78120
rect 207880 78100 208000 78120
rect 196000 78090 208000 78100
rect 196000 78020 196150 78090
rect 196350 78020 196650 78090
rect 196850 78020 197150 78090
rect 197350 78020 197650 78090
rect 197850 78020 198150 78090
rect 198350 78020 198650 78090
rect 198850 78020 199150 78090
rect 199350 78020 199650 78090
rect 199850 78020 200150 78090
rect 200350 78020 200650 78090
rect 200850 78020 201150 78090
rect 201350 78020 201650 78090
rect 201850 78020 202150 78090
rect 202350 78020 202650 78090
rect 202850 78020 203150 78090
rect 203350 78020 203650 78090
rect 203850 78020 204150 78090
rect 204350 78020 204650 78090
rect 204850 78020 205150 78090
rect 205350 78020 205650 78090
rect 205850 78020 206150 78090
rect 206350 78020 206650 78090
rect 206850 78020 207150 78090
rect 207350 78020 207650 78090
rect 207850 78020 208000 78090
rect 196000 77980 208000 78020
rect 196000 77910 196150 77980
rect 196350 77910 196650 77980
rect 196850 77910 197150 77980
rect 197350 77910 197650 77980
rect 197850 77910 198150 77980
rect 198350 77910 198650 77980
rect 198850 77910 199150 77980
rect 199350 77910 199650 77980
rect 199850 77910 200150 77980
rect 200350 77910 200650 77980
rect 200850 77910 201150 77980
rect 201350 77910 201650 77980
rect 201850 77910 202150 77980
rect 202350 77910 202650 77980
rect 202850 77910 203150 77980
rect 203350 77910 203650 77980
rect 203850 77910 204150 77980
rect 204350 77910 204650 77980
rect 204850 77910 205150 77980
rect 205350 77910 205650 77980
rect 205850 77910 206150 77980
rect 206350 77910 206650 77980
rect 206850 77910 207150 77980
rect 207350 77910 207650 77980
rect 207850 77910 208000 77980
rect 196000 77900 208000 77910
rect 196000 77880 196120 77900
rect 196380 77880 196620 77900
rect 196880 77880 197120 77900
rect 197380 77880 197620 77900
rect 197880 77880 198120 77900
rect 198380 77880 198620 77900
rect 198880 77880 199120 77900
rect 199380 77880 199620 77900
rect 199880 77880 200120 77900
rect 200380 77880 200620 77900
rect 200880 77880 201120 77900
rect 201380 77880 201620 77900
rect 201880 77880 202120 77900
rect 202380 77880 202620 77900
rect 202880 77880 203120 77900
rect 203380 77880 203620 77900
rect 203880 77880 204120 77900
rect 204380 77880 204620 77900
rect 204880 77880 205120 77900
rect 205380 77880 205620 77900
rect 205880 77880 206120 77900
rect 206380 77880 206620 77900
rect 206880 77880 207120 77900
rect 207380 77880 207620 77900
rect 207880 77880 208000 77900
rect 196000 77850 196100 77880
rect 196000 77650 196020 77850
rect 196090 77650 196100 77850
rect 196000 77620 196100 77650
rect 196400 77850 196600 77880
rect 196400 77650 196410 77850
rect 196480 77650 196520 77850
rect 196590 77650 196600 77850
rect 196400 77620 196600 77650
rect 196900 77850 197100 77880
rect 196900 77650 196910 77850
rect 196980 77650 197020 77850
rect 197090 77650 197100 77850
rect 196900 77620 197100 77650
rect 197400 77850 197600 77880
rect 197400 77650 197410 77850
rect 197480 77650 197520 77850
rect 197590 77650 197600 77850
rect 197400 77620 197600 77650
rect 197900 77850 198100 77880
rect 197900 77650 197910 77850
rect 197980 77650 198020 77850
rect 198090 77650 198100 77850
rect 197900 77620 198100 77650
rect 198400 77850 198600 77880
rect 198400 77650 198410 77850
rect 198480 77650 198520 77850
rect 198590 77650 198600 77850
rect 198400 77620 198600 77650
rect 198900 77850 199100 77880
rect 198900 77650 198910 77850
rect 198980 77650 199020 77850
rect 199090 77650 199100 77850
rect 198900 77620 199100 77650
rect 199400 77850 199600 77880
rect 199400 77650 199410 77850
rect 199480 77650 199520 77850
rect 199590 77650 199600 77850
rect 199400 77620 199600 77650
rect 199900 77850 200100 77880
rect 199900 77650 199910 77850
rect 199980 77650 200020 77850
rect 200090 77650 200100 77850
rect 199900 77620 200100 77650
rect 200400 77850 200600 77880
rect 200400 77650 200410 77850
rect 200480 77650 200520 77850
rect 200590 77650 200600 77850
rect 200400 77620 200600 77650
rect 200900 77850 201100 77880
rect 200900 77650 200910 77850
rect 200980 77650 201020 77850
rect 201090 77650 201100 77850
rect 200900 77620 201100 77650
rect 201400 77850 201600 77880
rect 201400 77650 201410 77850
rect 201480 77650 201520 77850
rect 201590 77650 201600 77850
rect 201400 77620 201600 77650
rect 201900 77850 202100 77880
rect 201900 77650 201910 77850
rect 201980 77650 202020 77850
rect 202090 77650 202100 77850
rect 201900 77620 202100 77650
rect 202400 77850 202600 77880
rect 202400 77650 202410 77850
rect 202480 77650 202520 77850
rect 202590 77650 202600 77850
rect 202400 77620 202600 77650
rect 202900 77850 203100 77880
rect 202900 77650 202910 77850
rect 202980 77650 203020 77850
rect 203090 77650 203100 77850
rect 202900 77620 203100 77650
rect 203400 77850 203600 77880
rect 203400 77650 203410 77850
rect 203480 77650 203520 77850
rect 203590 77650 203600 77850
rect 203400 77620 203600 77650
rect 203900 77850 204100 77880
rect 203900 77650 203910 77850
rect 203980 77650 204020 77850
rect 204090 77650 204100 77850
rect 203900 77620 204100 77650
rect 204400 77850 204600 77880
rect 204400 77650 204410 77850
rect 204480 77650 204520 77850
rect 204590 77650 204600 77850
rect 204400 77620 204600 77650
rect 204900 77850 205100 77880
rect 204900 77650 204910 77850
rect 204980 77650 205020 77850
rect 205090 77650 205100 77850
rect 204900 77620 205100 77650
rect 205400 77850 205600 77880
rect 205400 77650 205410 77850
rect 205480 77650 205520 77850
rect 205590 77650 205600 77850
rect 205400 77620 205600 77650
rect 205900 77850 206100 77880
rect 205900 77650 205910 77850
rect 205980 77650 206020 77850
rect 206090 77650 206100 77850
rect 205900 77620 206100 77650
rect 206400 77850 206600 77880
rect 206400 77650 206410 77850
rect 206480 77650 206520 77850
rect 206590 77650 206600 77850
rect 206400 77620 206600 77650
rect 206900 77850 207100 77880
rect 206900 77650 206910 77850
rect 206980 77650 207020 77850
rect 207090 77650 207100 77850
rect 206900 77620 207100 77650
rect 207400 77850 207600 77880
rect 207400 77650 207410 77850
rect 207480 77650 207520 77850
rect 207590 77650 207600 77850
rect 207400 77620 207600 77650
rect 207900 77850 208000 77880
rect 207900 77650 207910 77850
rect 207980 77650 208000 77850
rect 207900 77620 208000 77650
rect 196000 77600 196120 77620
rect 196380 77600 196620 77620
rect 196880 77600 197120 77620
rect 197380 77600 197620 77620
rect 197880 77600 198120 77620
rect 198380 77600 198620 77620
rect 198880 77600 199120 77620
rect 199380 77600 199620 77620
rect 199880 77600 200120 77620
rect 200380 77600 200620 77620
rect 200880 77600 201120 77620
rect 201380 77600 201620 77620
rect 201880 77600 202120 77620
rect 202380 77600 202620 77620
rect 202880 77600 203120 77620
rect 203380 77600 203620 77620
rect 203880 77600 204120 77620
rect 204380 77600 204620 77620
rect 204880 77600 205120 77620
rect 205380 77600 205620 77620
rect 205880 77600 206120 77620
rect 206380 77600 206620 77620
rect 206880 77600 207120 77620
rect 207380 77600 207620 77620
rect 207880 77600 208000 77620
rect 196000 77590 208000 77600
rect 196000 77520 196150 77590
rect 196350 77520 196650 77590
rect 196850 77520 197150 77590
rect 197350 77520 197650 77590
rect 197850 77520 198150 77590
rect 198350 77520 198650 77590
rect 198850 77520 199150 77590
rect 199350 77520 199650 77590
rect 199850 77520 200150 77590
rect 200350 77520 200650 77590
rect 200850 77520 201150 77590
rect 201350 77520 201650 77590
rect 201850 77520 202150 77590
rect 202350 77520 202650 77590
rect 202850 77520 203150 77590
rect 203350 77520 203650 77590
rect 203850 77520 204150 77590
rect 204350 77520 204650 77590
rect 204850 77520 205150 77590
rect 205350 77520 205650 77590
rect 205850 77520 206150 77590
rect 206350 77520 206650 77590
rect 206850 77520 207150 77590
rect 207350 77520 207650 77590
rect 207850 77520 208000 77590
rect 196000 77480 208000 77520
rect 196000 77410 196150 77480
rect 196350 77410 196650 77480
rect 196850 77410 197150 77480
rect 197350 77410 197650 77480
rect 197850 77410 198150 77480
rect 198350 77410 198650 77480
rect 198850 77410 199150 77480
rect 199350 77410 199650 77480
rect 199850 77410 200150 77480
rect 200350 77410 200650 77480
rect 200850 77410 201150 77480
rect 201350 77410 201650 77480
rect 201850 77410 202150 77480
rect 202350 77410 202650 77480
rect 202850 77410 203150 77480
rect 203350 77410 203650 77480
rect 203850 77410 204150 77480
rect 204350 77410 204650 77480
rect 204850 77410 205150 77480
rect 205350 77410 205650 77480
rect 205850 77410 206150 77480
rect 206350 77410 206650 77480
rect 206850 77410 207150 77480
rect 207350 77410 207650 77480
rect 207850 77410 208000 77480
rect 196000 77400 208000 77410
rect 196000 77380 196120 77400
rect 196380 77380 196620 77400
rect 196880 77380 197120 77400
rect 197380 77380 197620 77400
rect 197880 77380 198120 77400
rect 198380 77380 198620 77400
rect 198880 77380 199120 77400
rect 199380 77380 199620 77400
rect 199880 77380 200120 77400
rect 200380 77380 200620 77400
rect 200880 77380 201120 77400
rect 201380 77380 201620 77400
rect 201880 77380 202120 77400
rect 202380 77380 202620 77400
rect 202880 77380 203120 77400
rect 203380 77380 203620 77400
rect 203880 77380 204120 77400
rect 204380 77380 204620 77400
rect 204880 77380 205120 77400
rect 205380 77380 205620 77400
rect 205880 77380 206120 77400
rect 206380 77380 206620 77400
rect 206880 77380 207120 77400
rect 207380 77380 207620 77400
rect 207880 77380 208000 77400
rect 196000 77350 196100 77380
rect 196000 77150 196020 77350
rect 196090 77150 196100 77350
rect 196000 77120 196100 77150
rect 196400 77350 196600 77380
rect 196400 77150 196410 77350
rect 196480 77150 196520 77350
rect 196590 77150 196600 77350
rect 196400 77120 196600 77150
rect 196900 77350 197100 77380
rect 196900 77150 196910 77350
rect 196980 77150 197020 77350
rect 197090 77150 197100 77350
rect 196900 77120 197100 77150
rect 197400 77350 197600 77380
rect 197400 77150 197410 77350
rect 197480 77150 197520 77350
rect 197590 77150 197600 77350
rect 197400 77120 197600 77150
rect 197900 77350 198100 77380
rect 197900 77150 197910 77350
rect 197980 77150 198020 77350
rect 198090 77150 198100 77350
rect 197900 77120 198100 77150
rect 198400 77350 198600 77380
rect 198400 77150 198410 77350
rect 198480 77150 198520 77350
rect 198590 77150 198600 77350
rect 198400 77120 198600 77150
rect 198900 77350 199100 77380
rect 198900 77150 198910 77350
rect 198980 77150 199020 77350
rect 199090 77150 199100 77350
rect 198900 77120 199100 77150
rect 199400 77350 199600 77380
rect 199400 77150 199410 77350
rect 199480 77150 199520 77350
rect 199590 77150 199600 77350
rect 199400 77120 199600 77150
rect 199900 77350 200100 77380
rect 199900 77150 199910 77350
rect 199980 77150 200020 77350
rect 200090 77150 200100 77350
rect 199900 77120 200100 77150
rect 200400 77350 200600 77380
rect 200400 77150 200410 77350
rect 200480 77150 200520 77350
rect 200590 77150 200600 77350
rect 200400 77120 200600 77150
rect 200900 77350 201100 77380
rect 200900 77150 200910 77350
rect 200980 77150 201020 77350
rect 201090 77150 201100 77350
rect 200900 77120 201100 77150
rect 201400 77350 201600 77380
rect 201400 77150 201410 77350
rect 201480 77150 201520 77350
rect 201590 77150 201600 77350
rect 201400 77120 201600 77150
rect 201900 77350 202100 77380
rect 201900 77150 201910 77350
rect 201980 77150 202020 77350
rect 202090 77150 202100 77350
rect 201900 77120 202100 77150
rect 202400 77350 202600 77380
rect 202400 77150 202410 77350
rect 202480 77150 202520 77350
rect 202590 77150 202600 77350
rect 202400 77120 202600 77150
rect 202900 77350 203100 77380
rect 202900 77150 202910 77350
rect 202980 77150 203020 77350
rect 203090 77150 203100 77350
rect 202900 77120 203100 77150
rect 203400 77350 203600 77380
rect 203400 77150 203410 77350
rect 203480 77150 203520 77350
rect 203590 77150 203600 77350
rect 203400 77120 203600 77150
rect 203900 77350 204100 77380
rect 203900 77150 203910 77350
rect 203980 77150 204020 77350
rect 204090 77150 204100 77350
rect 203900 77120 204100 77150
rect 204400 77350 204600 77380
rect 204400 77150 204410 77350
rect 204480 77150 204520 77350
rect 204590 77150 204600 77350
rect 204400 77120 204600 77150
rect 204900 77350 205100 77380
rect 204900 77150 204910 77350
rect 204980 77150 205020 77350
rect 205090 77150 205100 77350
rect 204900 77120 205100 77150
rect 205400 77350 205600 77380
rect 205400 77150 205410 77350
rect 205480 77150 205520 77350
rect 205590 77150 205600 77350
rect 205400 77120 205600 77150
rect 205900 77350 206100 77380
rect 205900 77150 205910 77350
rect 205980 77150 206020 77350
rect 206090 77150 206100 77350
rect 205900 77120 206100 77150
rect 206400 77350 206600 77380
rect 206400 77150 206410 77350
rect 206480 77150 206520 77350
rect 206590 77150 206600 77350
rect 206400 77120 206600 77150
rect 206900 77350 207100 77380
rect 206900 77150 206910 77350
rect 206980 77150 207020 77350
rect 207090 77150 207100 77350
rect 206900 77120 207100 77150
rect 207400 77350 207600 77380
rect 207400 77150 207410 77350
rect 207480 77150 207520 77350
rect 207590 77150 207600 77350
rect 207400 77120 207600 77150
rect 207900 77350 208000 77380
rect 207900 77150 207910 77350
rect 207980 77150 208000 77350
rect 207900 77120 208000 77150
rect 196000 77100 196120 77120
rect 196380 77100 196620 77120
rect 196880 77100 197120 77120
rect 197380 77100 197620 77120
rect 197880 77100 198120 77120
rect 198380 77100 198620 77120
rect 198880 77100 199120 77120
rect 199380 77100 199620 77120
rect 199880 77100 200120 77120
rect 200380 77100 200620 77120
rect 200880 77100 201120 77120
rect 201380 77100 201620 77120
rect 201880 77100 202120 77120
rect 202380 77100 202620 77120
rect 202880 77100 203120 77120
rect 203380 77100 203620 77120
rect 203880 77100 204120 77120
rect 204380 77100 204620 77120
rect 204880 77100 205120 77120
rect 205380 77100 205620 77120
rect 205880 77100 206120 77120
rect 206380 77100 206620 77120
rect 206880 77100 207120 77120
rect 207380 77100 207620 77120
rect 207880 77100 208000 77120
rect 196000 77090 208000 77100
rect 196000 77020 196150 77090
rect 196350 77020 196650 77090
rect 196850 77020 197150 77090
rect 197350 77020 197650 77090
rect 197850 77020 198150 77090
rect 198350 77020 198650 77090
rect 198850 77020 199150 77090
rect 199350 77020 199650 77090
rect 199850 77020 200150 77090
rect 200350 77020 200650 77090
rect 200850 77020 201150 77090
rect 201350 77020 201650 77090
rect 201850 77020 202150 77090
rect 202350 77020 202650 77090
rect 202850 77020 203150 77090
rect 203350 77020 203650 77090
rect 203850 77020 204150 77090
rect 204350 77020 204650 77090
rect 204850 77020 205150 77090
rect 205350 77020 205650 77090
rect 205850 77020 206150 77090
rect 206350 77020 206650 77090
rect 206850 77020 207150 77090
rect 207350 77020 207650 77090
rect 207850 77020 208000 77090
rect 196000 76980 208000 77020
rect 196000 76910 196150 76980
rect 196350 76910 196650 76980
rect 196850 76910 197150 76980
rect 197350 76910 197650 76980
rect 197850 76910 198150 76980
rect 198350 76910 198650 76980
rect 198850 76910 199150 76980
rect 199350 76910 199650 76980
rect 199850 76910 200150 76980
rect 200350 76910 200650 76980
rect 200850 76910 201150 76980
rect 201350 76910 201650 76980
rect 201850 76910 202150 76980
rect 202350 76910 202650 76980
rect 202850 76910 203150 76980
rect 203350 76910 203650 76980
rect 203850 76910 204150 76980
rect 204350 76910 204650 76980
rect 204850 76910 205150 76980
rect 205350 76910 205650 76980
rect 205850 76910 206150 76980
rect 206350 76910 206650 76980
rect 206850 76910 207150 76980
rect 207350 76910 207650 76980
rect 207850 76910 208000 76980
rect 196000 76900 208000 76910
rect 196000 76880 196120 76900
rect 196380 76880 196620 76900
rect 196880 76880 197120 76900
rect 197380 76880 197620 76900
rect 197880 76880 198120 76900
rect 198380 76880 198620 76900
rect 198880 76880 199120 76900
rect 199380 76880 199620 76900
rect 199880 76880 200120 76900
rect 200380 76880 200620 76900
rect 200880 76880 201120 76900
rect 201380 76880 201620 76900
rect 201880 76880 202120 76900
rect 202380 76880 202620 76900
rect 202880 76880 203120 76900
rect 203380 76880 203620 76900
rect 203880 76880 204120 76900
rect 204380 76880 204620 76900
rect 204880 76880 205120 76900
rect 205380 76880 205620 76900
rect 205880 76880 206120 76900
rect 206380 76880 206620 76900
rect 206880 76880 207120 76900
rect 207380 76880 207620 76900
rect 207880 76880 208000 76900
rect 196000 76850 196100 76880
rect 196000 76650 196020 76850
rect 196090 76650 196100 76850
rect 196000 76620 196100 76650
rect 196400 76850 196600 76880
rect 196400 76650 196410 76850
rect 196480 76650 196520 76850
rect 196590 76650 196600 76850
rect 196400 76620 196600 76650
rect 196900 76850 197100 76880
rect 196900 76650 196910 76850
rect 196980 76650 197020 76850
rect 197090 76650 197100 76850
rect 196900 76620 197100 76650
rect 197400 76850 197600 76880
rect 197400 76650 197410 76850
rect 197480 76650 197520 76850
rect 197590 76650 197600 76850
rect 197400 76620 197600 76650
rect 197900 76850 198100 76880
rect 197900 76650 197910 76850
rect 197980 76650 198020 76850
rect 198090 76650 198100 76850
rect 197900 76620 198100 76650
rect 198400 76850 198600 76880
rect 198400 76650 198410 76850
rect 198480 76650 198520 76850
rect 198590 76650 198600 76850
rect 198400 76620 198600 76650
rect 198900 76850 199100 76880
rect 198900 76650 198910 76850
rect 198980 76650 199020 76850
rect 199090 76650 199100 76850
rect 198900 76620 199100 76650
rect 199400 76850 199600 76880
rect 199400 76650 199410 76850
rect 199480 76650 199520 76850
rect 199590 76650 199600 76850
rect 199400 76620 199600 76650
rect 199900 76850 200100 76880
rect 199900 76650 199910 76850
rect 199980 76650 200020 76850
rect 200090 76650 200100 76850
rect 199900 76620 200100 76650
rect 200400 76850 200600 76880
rect 200400 76650 200410 76850
rect 200480 76650 200520 76850
rect 200590 76650 200600 76850
rect 200400 76620 200600 76650
rect 200900 76850 201100 76880
rect 200900 76650 200910 76850
rect 200980 76650 201020 76850
rect 201090 76650 201100 76850
rect 200900 76620 201100 76650
rect 201400 76850 201600 76880
rect 201400 76650 201410 76850
rect 201480 76650 201520 76850
rect 201590 76650 201600 76850
rect 201400 76620 201600 76650
rect 201900 76850 202100 76880
rect 201900 76650 201910 76850
rect 201980 76650 202020 76850
rect 202090 76650 202100 76850
rect 201900 76620 202100 76650
rect 202400 76850 202600 76880
rect 202400 76650 202410 76850
rect 202480 76650 202520 76850
rect 202590 76650 202600 76850
rect 202400 76620 202600 76650
rect 202900 76850 203100 76880
rect 202900 76650 202910 76850
rect 202980 76650 203020 76850
rect 203090 76650 203100 76850
rect 202900 76620 203100 76650
rect 203400 76850 203600 76880
rect 203400 76650 203410 76850
rect 203480 76650 203520 76850
rect 203590 76650 203600 76850
rect 203400 76620 203600 76650
rect 203900 76850 204100 76880
rect 203900 76650 203910 76850
rect 203980 76650 204020 76850
rect 204090 76650 204100 76850
rect 203900 76620 204100 76650
rect 204400 76850 204600 76880
rect 204400 76650 204410 76850
rect 204480 76650 204520 76850
rect 204590 76650 204600 76850
rect 204400 76620 204600 76650
rect 204900 76850 205100 76880
rect 204900 76650 204910 76850
rect 204980 76650 205020 76850
rect 205090 76650 205100 76850
rect 204900 76620 205100 76650
rect 205400 76850 205600 76880
rect 205400 76650 205410 76850
rect 205480 76650 205520 76850
rect 205590 76650 205600 76850
rect 205400 76620 205600 76650
rect 205900 76850 206100 76880
rect 205900 76650 205910 76850
rect 205980 76650 206020 76850
rect 206090 76650 206100 76850
rect 205900 76620 206100 76650
rect 206400 76850 206600 76880
rect 206400 76650 206410 76850
rect 206480 76650 206520 76850
rect 206590 76650 206600 76850
rect 206400 76620 206600 76650
rect 206900 76850 207100 76880
rect 206900 76650 206910 76850
rect 206980 76650 207020 76850
rect 207090 76650 207100 76850
rect 206900 76620 207100 76650
rect 207400 76850 207600 76880
rect 207400 76650 207410 76850
rect 207480 76650 207520 76850
rect 207590 76650 207600 76850
rect 207400 76620 207600 76650
rect 207900 76850 208000 76880
rect 207900 76650 207910 76850
rect 207980 76650 208000 76850
rect 207900 76620 208000 76650
rect 196000 76600 196120 76620
rect 196380 76600 196620 76620
rect 196880 76600 197120 76620
rect 197380 76600 197620 76620
rect 197880 76600 198120 76620
rect 198380 76600 198620 76620
rect 198880 76600 199120 76620
rect 199380 76600 199620 76620
rect 199880 76600 200120 76620
rect 200380 76600 200620 76620
rect 200880 76600 201120 76620
rect 201380 76600 201620 76620
rect 201880 76600 202120 76620
rect 202380 76600 202620 76620
rect 202880 76600 203120 76620
rect 203380 76600 203620 76620
rect 203880 76600 204120 76620
rect 204380 76600 204620 76620
rect 204880 76600 205120 76620
rect 205380 76600 205620 76620
rect 205880 76600 206120 76620
rect 206380 76600 206620 76620
rect 206880 76600 207120 76620
rect 207380 76600 207620 76620
rect 207880 76600 208000 76620
rect 196000 76590 208000 76600
rect 196000 76520 196150 76590
rect 196350 76520 196650 76590
rect 196850 76520 197150 76590
rect 197350 76520 197650 76590
rect 197850 76520 198150 76590
rect 198350 76520 198650 76590
rect 198850 76520 199150 76590
rect 199350 76520 199650 76590
rect 199850 76520 200150 76590
rect 200350 76520 200650 76590
rect 200850 76520 201150 76590
rect 201350 76520 201650 76590
rect 201850 76520 202150 76590
rect 202350 76520 202650 76590
rect 202850 76520 203150 76590
rect 203350 76520 203650 76590
rect 203850 76520 204150 76590
rect 204350 76520 204650 76590
rect 204850 76520 205150 76590
rect 205350 76520 205650 76590
rect 205850 76520 206150 76590
rect 206350 76520 206650 76590
rect 206850 76520 207150 76590
rect 207350 76520 207650 76590
rect 207850 76520 208000 76590
rect 196000 76480 208000 76520
rect 196000 76410 196150 76480
rect 196350 76410 196650 76480
rect 196850 76410 197150 76480
rect 197350 76410 197650 76480
rect 197850 76410 198150 76480
rect 198350 76410 198650 76480
rect 198850 76410 199150 76480
rect 199350 76410 199650 76480
rect 199850 76410 200150 76480
rect 200350 76410 200650 76480
rect 200850 76410 201150 76480
rect 201350 76410 201650 76480
rect 201850 76410 202150 76480
rect 202350 76410 202650 76480
rect 202850 76410 203150 76480
rect 203350 76410 203650 76480
rect 203850 76410 204150 76480
rect 204350 76410 204650 76480
rect 204850 76410 205150 76480
rect 205350 76410 205650 76480
rect 205850 76410 206150 76480
rect 206350 76410 206650 76480
rect 206850 76410 207150 76480
rect 207350 76410 207650 76480
rect 207850 76410 208000 76480
rect 196000 76400 208000 76410
rect 196000 76380 196120 76400
rect 196380 76380 196620 76400
rect 196880 76380 197120 76400
rect 197380 76380 197620 76400
rect 197880 76380 198120 76400
rect 198380 76380 198620 76400
rect 198880 76380 199120 76400
rect 199380 76380 199620 76400
rect 199880 76380 200120 76400
rect 200380 76380 200620 76400
rect 200880 76380 201120 76400
rect 201380 76380 201620 76400
rect 201880 76380 202120 76400
rect 202380 76380 202620 76400
rect 202880 76380 203120 76400
rect 203380 76380 203620 76400
rect 203880 76380 204120 76400
rect 204380 76380 204620 76400
rect 204880 76380 205120 76400
rect 205380 76380 205620 76400
rect 205880 76380 206120 76400
rect 206380 76380 206620 76400
rect 206880 76380 207120 76400
rect 207380 76380 207620 76400
rect 207880 76380 208000 76400
rect 196000 76350 196100 76380
rect 196000 76150 196020 76350
rect 196090 76150 196100 76350
rect 196000 76120 196100 76150
rect 196400 76350 196600 76380
rect 196400 76150 196410 76350
rect 196480 76150 196520 76350
rect 196590 76150 196600 76350
rect 196400 76120 196600 76150
rect 196900 76350 197100 76380
rect 196900 76150 196910 76350
rect 196980 76150 197020 76350
rect 197090 76150 197100 76350
rect 196900 76120 197100 76150
rect 197400 76350 197600 76380
rect 197400 76150 197410 76350
rect 197480 76150 197520 76350
rect 197590 76150 197600 76350
rect 197400 76120 197600 76150
rect 197900 76350 198100 76380
rect 197900 76150 197910 76350
rect 197980 76150 198020 76350
rect 198090 76150 198100 76350
rect 197900 76120 198100 76150
rect 198400 76350 198600 76380
rect 198400 76150 198410 76350
rect 198480 76150 198520 76350
rect 198590 76150 198600 76350
rect 198400 76120 198600 76150
rect 198900 76350 199100 76380
rect 198900 76150 198910 76350
rect 198980 76150 199020 76350
rect 199090 76150 199100 76350
rect 198900 76120 199100 76150
rect 199400 76350 199600 76380
rect 199400 76150 199410 76350
rect 199480 76150 199520 76350
rect 199590 76150 199600 76350
rect 199400 76120 199600 76150
rect 199900 76350 200100 76380
rect 199900 76150 199910 76350
rect 199980 76150 200020 76350
rect 200090 76150 200100 76350
rect 199900 76120 200100 76150
rect 200400 76350 200600 76380
rect 200400 76150 200410 76350
rect 200480 76150 200520 76350
rect 200590 76150 200600 76350
rect 200400 76120 200600 76150
rect 200900 76350 201100 76380
rect 200900 76150 200910 76350
rect 200980 76150 201020 76350
rect 201090 76150 201100 76350
rect 200900 76120 201100 76150
rect 201400 76350 201600 76380
rect 201400 76150 201410 76350
rect 201480 76150 201520 76350
rect 201590 76150 201600 76350
rect 201400 76120 201600 76150
rect 201900 76350 202100 76380
rect 201900 76150 201910 76350
rect 201980 76150 202020 76350
rect 202090 76150 202100 76350
rect 201900 76120 202100 76150
rect 202400 76350 202600 76380
rect 202400 76150 202410 76350
rect 202480 76150 202520 76350
rect 202590 76150 202600 76350
rect 202400 76120 202600 76150
rect 202900 76350 203100 76380
rect 202900 76150 202910 76350
rect 202980 76150 203020 76350
rect 203090 76150 203100 76350
rect 202900 76120 203100 76150
rect 203400 76350 203600 76380
rect 203400 76150 203410 76350
rect 203480 76150 203520 76350
rect 203590 76150 203600 76350
rect 203400 76120 203600 76150
rect 203900 76350 204100 76380
rect 203900 76150 203910 76350
rect 203980 76150 204020 76350
rect 204090 76150 204100 76350
rect 203900 76120 204100 76150
rect 204400 76350 204600 76380
rect 204400 76150 204410 76350
rect 204480 76150 204520 76350
rect 204590 76150 204600 76350
rect 204400 76120 204600 76150
rect 204900 76350 205100 76380
rect 204900 76150 204910 76350
rect 204980 76150 205020 76350
rect 205090 76150 205100 76350
rect 204900 76120 205100 76150
rect 205400 76350 205600 76380
rect 205400 76150 205410 76350
rect 205480 76150 205520 76350
rect 205590 76150 205600 76350
rect 205400 76120 205600 76150
rect 205900 76350 206100 76380
rect 205900 76150 205910 76350
rect 205980 76150 206020 76350
rect 206090 76150 206100 76350
rect 205900 76120 206100 76150
rect 206400 76350 206600 76380
rect 206400 76150 206410 76350
rect 206480 76150 206520 76350
rect 206590 76150 206600 76350
rect 206400 76120 206600 76150
rect 206900 76350 207100 76380
rect 206900 76150 206910 76350
rect 206980 76150 207020 76350
rect 207090 76150 207100 76350
rect 206900 76120 207100 76150
rect 207400 76350 207600 76380
rect 207400 76150 207410 76350
rect 207480 76150 207520 76350
rect 207590 76150 207600 76350
rect 207400 76120 207600 76150
rect 207900 76350 208000 76380
rect 207900 76150 207910 76350
rect 207980 76150 208000 76350
rect 207900 76120 208000 76150
rect 196000 76100 196120 76120
rect 196380 76100 196620 76120
rect 196880 76100 197120 76120
rect 197380 76100 197620 76120
rect 197880 76100 198120 76120
rect 198380 76100 198620 76120
rect 198880 76100 199120 76120
rect 199380 76100 199620 76120
rect 199880 76100 200120 76120
rect 200380 76100 200620 76120
rect 200880 76100 201120 76120
rect 201380 76100 201620 76120
rect 201880 76100 202120 76120
rect 202380 76100 202620 76120
rect 202880 76100 203120 76120
rect 203380 76100 203620 76120
rect 203880 76100 204120 76120
rect 204380 76100 204620 76120
rect 204880 76100 205120 76120
rect 205380 76100 205620 76120
rect 205880 76100 206120 76120
rect 206380 76100 206620 76120
rect 206880 76100 207120 76120
rect 207380 76100 207620 76120
rect 207880 76100 208000 76120
rect 196000 76090 208000 76100
rect 196000 76020 196150 76090
rect 196350 76020 196650 76090
rect 196850 76020 197150 76090
rect 197350 76020 197650 76090
rect 197850 76020 198150 76090
rect 198350 76020 198650 76090
rect 198850 76020 199150 76090
rect 199350 76020 199650 76090
rect 199850 76020 200150 76090
rect 200350 76020 200650 76090
rect 200850 76020 201150 76090
rect 201350 76020 201650 76090
rect 201850 76020 202150 76090
rect 202350 76020 202650 76090
rect 202850 76020 203150 76090
rect 203350 76020 203650 76090
rect 203850 76020 204150 76090
rect 204350 76020 204650 76090
rect 204850 76020 205150 76090
rect 205350 76020 205650 76090
rect 205850 76020 206150 76090
rect 206350 76020 206650 76090
rect 206850 76020 207150 76090
rect 207350 76020 207650 76090
rect 207850 76020 208000 76090
rect 196000 75980 208000 76020
rect 196000 75910 196150 75980
rect 196350 75910 196650 75980
rect 196850 75910 197150 75980
rect 197350 75910 197650 75980
rect 197850 75910 198150 75980
rect 198350 75910 198650 75980
rect 198850 75910 199150 75980
rect 199350 75910 199650 75980
rect 199850 75910 200150 75980
rect 200350 75910 200650 75980
rect 200850 75910 201150 75980
rect 201350 75910 201650 75980
rect 201850 75910 202150 75980
rect 202350 75910 202650 75980
rect 202850 75910 203150 75980
rect 203350 75910 203650 75980
rect 203850 75910 204150 75980
rect 204350 75910 204650 75980
rect 204850 75910 205150 75980
rect 205350 75910 205650 75980
rect 205850 75910 206150 75980
rect 206350 75910 206650 75980
rect 206850 75910 207150 75980
rect 207350 75910 207650 75980
rect 207850 75910 208000 75980
rect 196000 75900 208000 75910
rect 196000 75880 196120 75900
rect 196380 75880 196620 75900
rect 196880 75880 197120 75900
rect 197380 75880 197620 75900
rect 197880 75880 198120 75900
rect 198380 75880 198620 75900
rect 198880 75880 199120 75900
rect 199380 75880 199620 75900
rect 199880 75880 200120 75900
rect 200380 75880 200620 75900
rect 200880 75880 201120 75900
rect 201380 75880 201620 75900
rect 201880 75880 202120 75900
rect 202380 75880 202620 75900
rect 202880 75880 203120 75900
rect 203380 75880 203620 75900
rect 203880 75880 204120 75900
rect 204380 75880 204620 75900
rect 204880 75880 205120 75900
rect 205380 75880 205620 75900
rect 205880 75880 206120 75900
rect 206380 75880 206620 75900
rect 206880 75880 207120 75900
rect 207380 75880 207620 75900
rect 207880 75880 208000 75900
rect 196000 75850 196100 75880
rect 196000 75650 196020 75850
rect 196090 75650 196100 75850
rect 196000 75620 196100 75650
rect 196400 75850 196600 75880
rect 196400 75650 196410 75850
rect 196480 75650 196520 75850
rect 196590 75650 196600 75850
rect 196400 75620 196600 75650
rect 196900 75850 197100 75880
rect 196900 75650 196910 75850
rect 196980 75650 197020 75850
rect 197090 75650 197100 75850
rect 196900 75620 197100 75650
rect 197400 75850 197600 75880
rect 197400 75650 197410 75850
rect 197480 75650 197520 75850
rect 197590 75650 197600 75850
rect 197400 75620 197600 75650
rect 197900 75850 198100 75880
rect 197900 75650 197910 75850
rect 197980 75650 198020 75850
rect 198090 75650 198100 75850
rect 197900 75620 198100 75650
rect 198400 75850 198600 75880
rect 198400 75650 198410 75850
rect 198480 75650 198520 75850
rect 198590 75650 198600 75850
rect 198400 75620 198600 75650
rect 198900 75850 199100 75880
rect 198900 75650 198910 75850
rect 198980 75650 199020 75850
rect 199090 75650 199100 75850
rect 198900 75620 199100 75650
rect 199400 75850 199600 75880
rect 199400 75650 199410 75850
rect 199480 75650 199520 75850
rect 199590 75650 199600 75850
rect 199400 75620 199600 75650
rect 199900 75850 200100 75880
rect 199900 75650 199910 75850
rect 199980 75650 200020 75850
rect 200090 75650 200100 75850
rect 199900 75620 200100 75650
rect 200400 75850 200600 75880
rect 200400 75650 200410 75850
rect 200480 75650 200520 75850
rect 200590 75650 200600 75850
rect 200400 75620 200600 75650
rect 200900 75850 201100 75880
rect 200900 75650 200910 75850
rect 200980 75650 201020 75850
rect 201090 75650 201100 75850
rect 200900 75620 201100 75650
rect 201400 75850 201600 75880
rect 201400 75650 201410 75850
rect 201480 75650 201520 75850
rect 201590 75650 201600 75850
rect 201400 75620 201600 75650
rect 201900 75850 202100 75880
rect 201900 75650 201910 75850
rect 201980 75650 202020 75850
rect 202090 75650 202100 75850
rect 201900 75620 202100 75650
rect 202400 75850 202600 75880
rect 202400 75650 202410 75850
rect 202480 75650 202520 75850
rect 202590 75650 202600 75850
rect 202400 75620 202600 75650
rect 202900 75850 203100 75880
rect 202900 75650 202910 75850
rect 202980 75650 203020 75850
rect 203090 75650 203100 75850
rect 202900 75620 203100 75650
rect 203400 75850 203600 75880
rect 203400 75650 203410 75850
rect 203480 75650 203520 75850
rect 203590 75650 203600 75850
rect 203400 75620 203600 75650
rect 203900 75850 204100 75880
rect 203900 75650 203910 75850
rect 203980 75650 204020 75850
rect 204090 75650 204100 75850
rect 203900 75620 204100 75650
rect 204400 75850 204600 75880
rect 204400 75650 204410 75850
rect 204480 75650 204520 75850
rect 204590 75650 204600 75850
rect 204400 75620 204600 75650
rect 204900 75850 205100 75880
rect 204900 75650 204910 75850
rect 204980 75650 205020 75850
rect 205090 75650 205100 75850
rect 204900 75620 205100 75650
rect 205400 75850 205600 75880
rect 205400 75650 205410 75850
rect 205480 75650 205520 75850
rect 205590 75650 205600 75850
rect 205400 75620 205600 75650
rect 205900 75850 206100 75880
rect 205900 75650 205910 75850
rect 205980 75650 206020 75850
rect 206090 75650 206100 75850
rect 205900 75620 206100 75650
rect 206400 75850 206600 75880
rect 206400 75650 206410 75850
rect 206480 75650 206520 75850
rect 206590 75650 206600 75850
rect 206400 75620 206600 75650
rect 206900 75850 207100 75880
rect 206900 75650 206910 75850
rect 206980 75650 207020 75850
rect 207090 75650 207100 75850
rect 206900 75620 207100 75650
rect 207400 75850 207600 75880
rect 207400 75650 207410 75850
rect 207480 75650 207520 75850
rect 207590 75650 207600 75850
rect 207400 75620 207600 75650
rect 207900 75850 208000 75880
rect 207900 75650 207910 75850
rect 207980 75650 208000 75850
rect 207900 75620 208000 75650
rect 196000 75600 196120 75620
rect 196380 75600 196620 75620
rect 196880 75600 197120 75620
rect 197380 75600 197620 75620
rect 197880 75600 198120 75620
rect 198380 75600 198620 75620
rect 198880 75600 199120 75620
rect 199380 75600 199620 75620
rect 199880 75600 200120 75620
rect 200380 75600 200620 75620
rect 200880 75600 201120 75620
rect 201380 75600 201620 75620
rect 201880 75600 202120 75620
rect 202380 75600 202620 75620
rect 202880 75600 203120 75620
rect 203380 75600 203620 75620
rect 203880 75600 204120 75620
rect 204380 75600 204620 75620
rect 204880 75600 205120 75620
rect 205380 75600 205620 75620
rect 205880 75600 206120 75620
rect 206380 75600 206620 75620
rect 206880 75600 207120 75620
rect 207380 75600 207620 75620
rect 207880 75600 208000 75620
rect 196000 75590 208000 75600
rect 196000 75520 196150 75590
rect 196350 75520 196650 75590
rect 196850 75520 197150 75590
rect 197350 75520 197650 75590
rect 197850 75520 198150 75590
rect 198350 75520 198650 75590
rect 198850 75520 199150 75590
rect 199350 75520 199650 75590
rect 199850 75520 200150 75590
rect 200350 75520 200650 75590
rect 200850 75520 201150 75590
rect 201350 75520 201650 75590
rect 201850 75520 202150 75590
rect 202350 75520 202650 75590
rect 202850 75520 203150 75590
rect 203350 75520 203650 75590
rect 203850 75520 204150 75590
rect 204350 75520 204650 75590
rect 204850 75520 205150 75590
rect 205350 75520 205650 75590
rect 205850 75520 206150 75590
rect 206350 75520 206650 75590
rect 206850 75520 207150 75590
rect 207350 75520 207650 75590
rect 207850 75520 208000 75590
rect 196000 75480 208000 75520
rect 196000 75410 196150 75480
rect 196350 75410 196650 75480
rect 196850 75410 197150 75480
rect 197350 75410 197650 75480
rect 197850 75410 198150 75480
rect 198350 75410 198650 75480
rect 198850 75410 199150 75480
rect 199350 75410 199650 75480
rect 199850 75410 200150 75480
rect 200350 75410 200650 75480
rect 200850 75410 201150 75480
rect 201350 75410 201650 75480
rect 201850 75410 202150 75480
rect 202350 75410 202650 75480
rect 202850 75410 203150 75480
rect 203350 75410 203650 75480
rect 203850 75410 204150 75480
rect 204350 75410 204650 75480
rect 204850 75410 205150 75480
rect 205350 75410 205650 75480
rect 205850 75410 206150 75480
rect 206350 75410 206650 75480
rect 206850 75410 207150 75480
rect 207350 75410 207650 75480
rect 207850 75410 208000 75480
rect 196000 75400 208000 75410
rect 196000 75380 196120 75400
rect 196380 75380 196620 75400
rect 196880 75380 197120 75400
rect 197380 75380 197620 75400
rect 197880 75380 198120 75400
rect 198380 75380 198620 75400
rect 198880 75380 199120 75400
rect 199380 75380 199620 75400
rect 199880 75380 200120 75400
rect 200380 75380 200620 75400
rect 200880 75380 201120 75400
rect 201380 75380 201620 75400
rect 201880 75380 202120 75400
rect 202380 75380 202620 75400
rect 202880 75380 203120 75400
rect 203380 75380 203620 75400
rect 203880 75380 204120 75400
rect 204380 75380 204620 75400
rect 204880 75380 205120 75400
rect 205380 75380 205620 75400
rect 205880 75380 206120 75400
rect 206380 75380 206620 75400
rect 206880 75380 207120 75400
rect 207380 75380 207620 75400
rect 207880 75380 208000 75400
rect 196000 75350 196100 75380
rect 196000 75150 196020 75350
rect 196090 75150 196100 75350
rect 196000 75120 196100 75150
rect 196400 75350 196600 75380
rect 196400 75150 196410 75350
rect 196480 75150 196520 75350
rect 196590 75150 196600 75350
rect 196400 75120 196600 75150
rect 196900 75350 197100 75380
rect 196900 75150 196910 75350
rect 196980 75150 197020 75350
rect 197090 75150 197100 75350
rect 196900 75120 197100 75150
rect 197400 75350 197600 75380
rect 197400 75150 197410 75350
rect 197480 75150 197520 75350
rect 197590 75150 197600 75350
rect 197400 75120 197600 75150
rect 197900 75350 198100 75380
rect 197900 75150 197910 75350
rect 197980 75150 198020 75350
rect 198090 75150 198100 75350
rect 197900 75120 198100 75150
rect 198400 75350 198600 75380
rect 198400 75150 198410 75350
rect 198480 75150 198520 75350
rect 198590 75150 198600 75350
rect 198400 75120 198600 75150
rect 198900 75350 199100 75380
rect 198900 75150 198910 75350
rect 198980 75150 199020 75350
rect 199090 75150 199100 75350
rect 198900 75120 199100 75150
rect 199400 75350 199600 75380
rect 199400 75150 199410 75350
rect 199480 75150 199520 75350
rect 199590 75150 199600 75350
rect 199400 75120 199600 75150
rect 199900 75350 200100 75380
rect 199900 75150 199910 75350
rect 199980 75150 200020 75350
rect 200090 75150 200100 75350
rect 199900 75120 200100 75150
rect 200400 75350 200600 75380
rect 200400 75150 200410 75350
rect 200480 75150 200520 75350
rect 200590 75150 200600 75350
rect 200400 75120 200600 75150
rect 200900 75350 201100 75380
rect 200900 75150 200910 75350
rect 200980 75150 201020 75350
rect 201090 75150 201100 75350
rect 200900 75120 201100 75150
rect 201400 75350 201600 75380
rect 201400 75150 201410 75350
rect 201480 75150 201520 75350
rect 201590 75150 201600 75350
rect 201400 75120 201600 75150
rect 201900 75350 202100 75380
rect 201900 75150 201910 75350
rect 201980 75150 202020 75350
rect 202090 75150 202100 75350
rect 201900 75120 202100 75150
rect 202400 75350 202600 75380
rect 202400 75150 202410 75350
rect 202480 75150 202520 75350
rect 202590 75150 202600 75350
rect 202400 75120 202600 75150
rect 202900 75350 203100 75380
rect 202900 75150 202910 75350
rect 202980 75150 203020 75350
rect 203090 75150 203100 75350
rect 202900 75120 203100 75150
rect 203400 75350 203600 75380
rect 203400 75150 203410 75350
rect 203480 75150 203520 75350
rect 203590 75150 203600 75350
rect 203400 75120 203600 75150
rect 203900 75350 204100 75380
rect 203900 75150 203910 75350
rect 203980 75150 204020 75350
rect 204090 75150 204100 75350
rect 203900 75120 204100 75150
rect 204400 75350 204600 75380
rect 204400 75150 204410 75350
rect 204480 75150 204520 75350
rect 204590 75150 204600 75350
rect 204400 75120 204600 75150
rect 204900 75350 205100 75380
rect 204900 75150 204910 75350
rect 204980 75150 205020 75350
rect 205090 75150 205100 75350
rect 204900 75120 205100 75150
rect 205400 75350 205600 75380
rect 205400 75150 205410 75350
rect 205480 75150 205520 75350
rect 205590 75150 205600 75350
rect 205400 75120 205600 75150
rect 205900 75350 206100 75380
rect 205900 75150 205910 75350
rect 205980 75150 206020 75350
rect 206090 75150 206100 75350
rect 205900 75120 206100 75150
rect 206400 75350 206600 75380
rect 206400 75150 206410 75350
rect 206480 75150 206520 75350
rect 206590 75150 206600 75350
rect 206400 75120 206600 75150
rect 206900 75350 207100 75380
rect 206900 75150 206910 75350
rect 206980 75150 207020 75350
rect 207090 75150 207100 75350
rect 206900 75120 207100 75150
rect 207400 75350 207600 75380
rect 207400 75150 207410 75350
rect 207480 75150 207520 75350
rect 207590 75150 207600 75350
rect 207400 75120 207600 75150
rect 207900 75350 208000 75380
rect 207900 75150 207910 75350
rect 207980 75150 208000 75350
rect 207900 75120 208000 75150
rect 196000 75100 196120 75120
rect 196380 75100 196620 75120
rect 196880 75100 197120 75120
rect 197380 75100 197620 75120
rect 197880 75100 198120 75120
rect 198380 75100 198620 75120
rect 198880 75100 199120 75120
rect 199380 75100 199620 75120
rect 199880 75100 200120 75120
rect 200380 75100 200620 75120
rect 200880 75100 201120 75120
rect 201380 75100 201620 75120
rect 201880 75100 202120 75120
rect 202380 75100 202620 75120
rect 202880 75100 203120 75120
rect 203380 75100 203620 75120
rect 203880 75100 204120 75120
rect 204380 75100 204620 75120
rect 204880 75100 205120 75120
rect 205380 75100 205620 75120
rect 205880 75100 206120 75120
rect 206380 75100 206620 75120
rect 206880 75100 207120 75120
rect 207380 75100 207620 75120
rect 207880 75100 208000 75120
rect 196000 75090 208000 75100
rect 196000 75020 196150 75090
rect 196350 75020 196650 75090
rect 196850 75020 197150 75090
rect 197350 75020 197650 75090
rect 197850 75020 198150 75090
rect 198350 75020 198650 75090
rect 198850 75020 199150 75090
rect 199350 75020 199650 75090
rect 199850 75020 200150 75090
rect 200350 75020 200650 75090
rect 200850 75020 201150 75090
rect 201350 75020 201650 75090
rect 201850 75020 202150 75090
rect 202350 75020 202650 75090
rect 202850 75020 203150 75090
rect 203350 75020 203650 75090
rect 203850 75020 204150 75090
rect 204350 75020 204650 75090
rect 204850 75020 205150 75090
rect 205350 75020 205650 75090
rect 205850 75020 206150 75090
rect 206350 75020 206650 75090
rect 206850 75020 207150 75090
rect 207350 75020 207650 75090
rect 207850 75020 208000 75090
rect 196000 74980 208000 75020
rect 196000 74910 196150 74980
rect 196350 74910 196650 74980
rect 196850 74910 197150 74980
rect 197350 74910 197650 74980
rect 197850 74910 198150 74980
rect 198350 74910 198650 74980
rect 198850 74910 199150 74980
rect 199350 74910 199650 74980
rect 199850 74910 200150 74980
rect 200350 74910 200650 74980
rect 200850 74910 201150 74980
rect 201350 74910 201650 74980
rect 201850 74910 202150 74980
rect 202350 74910 202650 74980
rect 202850 74910 203150 74980
rect 203350 74910 203650 74980
rect 203850 74910 204150 74980
rect 204350 74910 204650 74980
rect 204850 74910 205150 74980
rect 205350 74910 205650 74980
rect 205850 74910 206150 74980
rect 206350 74910 206650 74980
rect 206850 74910 207150 74980
rect 207350 74910 207650 74980
rect 207850 74910 208000 74980
rect 196000 74900 208000 74910
rect 196000 74880 196120 74900
rect 196380 74880 196620 74900
rect 196880 74880 197120 74900
rect 197380 74880 197620 74900
rect 197880 74880 198120 74900
rect 198380 74880 198620 74900
rect 198880 74880 199120 74900
rect 199380 74880 199620 74900
rect 199880 74880 200120 74900
rect 200380 74880 200620 74900
rect 200880 74880 201120 74900
rect 201380 74880 201620 74900
rect 201880 74880 202120 74900
rect 202380 74880 202620 74900
rect 202880 74880 203120 74900
rect 203380 74880 203620 74900
rect 203880 74880 204120 74900
rect 204380 74880 204620 74900
rect 204880 74880 205120 74900
rect 205380 74880 205620 74900
rect 205880 74880 206120 74900
rect 206380 74880 206620 74900
rect 206880 74880 207120 74900
rect 207380 74880 207620 74900
rect 207880 74880 208000 74900
rect 196000 74850 196100 74880
rect 196000 74650 196020 74850
rect 196090 74650 196100 74850
rect 196000 74620 196100 74650
rect 196400 74850 196600 74880
rect 196400 74650 196410 74850
rect 196480 74650 196520 74850
rect 196590 74650 196600 74850
rect 196400 74620 196600 74650
rect 196900 74850 197100 74880
rect 196900 74650 196910 74850
rect 196980 74650 197020 74850
rect 197090 74650 197100 74850
rect 196900 74620 197100 74650
rect 197400 74850 197600 74880
rect 197400 74650 197410 74850
rect 197480 74650 197520 74850
rect 197590 74650 197600 74850
rect 197400 74620 197600 74650
rect 197900 74850 198100 74880
rect 197900 74650 197910 74850
rect 197980 74650 198020 74850
rect 198090 74650 198100 74850
rect 197900 74620 198100 74650
rect 198400 74850 198600 74880
rect 198400 74650 198410 74850
rect 198480 74650 198520 74850
rect 198590 74650 198600 74850
rect 198400 74620 198600 74650
rect 198900 74850 199100 74880
rect 198900 74650 198910 74850
rect 198980 74650 199020 74850
rect 199090 74650 199100 74850
rect 198900 74620 199100 74650
rect 199400 74850 199600 74880
rect 199400 74650 199410 74850
rect 199480 74650 199520 74850
rect 199590 74650 199600 74850
rect 199400 74620 199600 74650
rect 199900 74850 200100 74880
rect 199900 74650 199910 74850
rect 199980 74650 200020 74850
rect 200090 74650 200100 74850
rect 199900 74620 200100 74650
rect 200400 74850 200600 74880
rect 200400 74650 200410 74850
rect 200480 74650 200520 74850
rect 200590 74650 200600 74850
rect 200400 74620 200600 74650
rect 200900 74850 201100 74880
rect 200900 74650 200910 74850
rect 200980 74650 201020 74850
rect 201090 74650 201100 74850
rect 200900 74620 201100 74650
rect 201400 74850 201600 74880
rect 201400 74650 201410 74850
rect 201480 74650 201520 74850
rect 201590 74650 201600 74850
rect 201400 74620 201600 74650
rect 201900 74850 202100 74880
rect 201900 74650 201910 74850
rect 201980 74650 202020 74850
rect 202090 74650 202100 74850
rect 201900 74620 202100 74650
rect 202400 74850 202600 74880
rect 202400 74650 202410 74850
rect 202480 74650 202520 74850
rect 202590 74650 202600 74850
rect 202400 74620 202600 74650
rect 202900 74850 203100 74880
rect 202900 74650 202910 74850
rect 202980 74650 203020 74850
rect 203090 74650 203100 74850
rect 202900 74620 203100 74650
rect 203400 74850 203600 74880
rect 203400 74650 203410 74850
rect 203480 74650 203520 74850
rect 203590 74650 203600 74850
rect 203400 74620 203600 74650
rect 203900 74850 204100 74880
rect 203900 74650 203910 74850
rect 203980 74650 204020 74850
rect 204090 74650 204100 74850
rect 203900 74620 204100 74650
rect 204400 74850 204600 74880
rect 204400 74650 204410 74850
rect 204480 74650 204520 74850
rect 204590 74650 204600 74850
rect 204400 74620 204600 74650
rect 204900 74850 205100 74880
rect 204900 74650 204910 74850
rect 204980 74650 205020 74850
rect 205090 74650 205100 74850
rect 204900 74620 205100 74650
rect 205400 74850 205600 74880
rect 205400 74650 205410 74850
rect 205480 74650 205520 74850
rect 205590 74650 205600 74850
rect 205400 74620 205600 74650
rect 205900 74850 206100 74880
rect 205900 74650 205910 74850
rect 205980 74650 206020 74850
rect 206090 74650 206100 74850
rect 205900 74620 206100 74650
rect 206400 74850 206600 74880
rect 206400 74650 206410 74850
rect 206480 74650 206520 74850
rect 206590 74650 206600 74850
rect 206400 74620 206600 74650
rect 206900 74850 207100 74880
rect 206900 74650 206910 74850
rect 206980 74650 207020 74850
rect 207090 74650 207100 74850
rect 206900 74620 207100 74650
rect 207400 74850 207600 74880
rect 207400 74650 207410 74850
rect 207480 74650 207520 74850
rect 207590 74650 207600 74850
rect 207400 74620 207600 74650
rect 207900 74850 208000 74880
rect 207900 74650 207910 74850
rect 207980 74650 208000 74850
rect 207900 74620 208000 74650
rect 196000 74600 196120 74620
rect 196380 74600 196620 74620
rect 196880 74600 197120 74620
rect 197380 74600 197620 74620
rect 197880 74600 198120 74620
rect 198380 74600 198620 74620
rect 198880 74600 199120 74620
rect 199380 74600 199620 74620
rect 199880 74600 200120 74620
rect 200380 74600 200620 74620
rect 200880 74600 201120 74620
rect 201380 74600 201620 74620
rect 201880 74600 202120 74620
rect 202380 74600 202620 74620
rect 202880 74600 203120 74620
rect 203380 74600 203620 74620
rect 203880 74600 204120 74620
rect 204380 74600 204620 74620
rect 204880 74600 205120 74620
rect 205380 74600 205620 74620
rect 205880 74600 206120 74620
rect 206380 74600 206620 74620
rect 206880 74600 207120 74620
rect 207380 74600 207620 74620
rect 207880 74600 208000 74620
rect 196000 74590 208000 74600
rect 196000 74520 196150 74590
rect 196350 74520 196650 74590
rect 196850 74520 197150 74590
rect 197350 74520 197650 74590
rect 197850 74520 198150 74590
rect 198350 74520 198650 74590
rect 198850 74520 199150 74590
rect 199350 74520 199650 74590
rect 199850 74520 200150 74590
rect 200350 74520 200650 74590
rect 200850 74520 201150 74590
rect 201350 74520 201650 74590
rect 201850 74520 202150 74590
rect 202350 74520 202650 74590
rect 202850 74520 203150 74590
rect 203350 74520 203650 74590
rect 203850 74520 204150 74590
rect 204350 74520 204650 74590
rect 204850 74520 205150 74590
rect 205350 74520 205650 74590
rect 205850 74520 206150 74590
rect 206350 74520 206650 74590
rect 206850 74520 207150 74590
rect 207350 74520 207650 74590
rect 207850 74520 208000 74590
rect 196000 74480 208000 74520
rect 196000 74410 196150 74480
rect 196350 74410 196650 74480
rect 196850 74410 197150 74480
rect 197350 74410 197650 74480
rect 197850 74410 198150 74480
rect 198350 74410 198650 74480
rect 198850 74410 199150 74480
rect 199350 74410 199650 74480
rect 199850 74410 200150 74480
rect 200350 74410 200650 74480
rect 200850 74410 201150 74480
rect 201350 74410 201650 74480
rect 201850 74410 202150 74480
rect 202350 74410 202650 74480
rect 202850 74410 203150 74480
rect 203350 74410 203650 74480
rect 203850 74410 204150 74480
rect 204350 74410 204650 74480
rect 204850 74410 205150 74480
rect 205350 74410 205650 74480
rect 205850 74410 206150 74480
rect 206350 74410 206650 74480
rect 206850 74410 207150 74480
rect 207350 74410 207650 74480
rect 207850 74410 208000 74480
rect 196000 74400 208000 74410
rect 196000 74380 196120 74400
rect 196380 74380 196620 74400
rect 196880 74380 197120 74400
rect 197380 74380 197620 74400
rect 197880 74380 198120 74400
rect 198380 74380 198620 74400
rect 198880 74380 199120 74400
rect 199380 74380 199620 74400
rect 199880 74380 200120 74400
rect 200380 74380 200620 74400
rect 200880 74380 201120 74400
rect 201380 74380 201620 74400
rect 201880 74380 202120 74400
rect 202380 74380 202620 74400
rect 202880 74380 203120 74400
rect 203380 74380 203620 74400
rect 203880 74380 204120 74400
rect 204380 74380 204620 74400
rect 204880 74380 205120 74400
rect 205380 74380 205620 74400
rect 205880 74380 206120 74400
rect 206380 74380 206620 74400
rect 206880 74380 207120 74400
rect 207380 74380 207620 74400
rect 207880 74380 208000 74400
rect 196000 74350 196100 74380
rect 196000 74150 196020 74350
rect 196090 74150 196100 74350
rect 196000 74120 196100 74150
rect 196400 74350 196600 74380
rect 196400 74150 196410 74350
rect 196480 74150 196520 74350
rect 196590 74150 196600 74350
rect 196400 74120 196600 74150
rect 196900 74350 197100 74380
rect 196900 74150 196910 74350
rect 196980 74150 197020 74350
rect 197090 74150 197100 74350
rect 196900 74120 197100 74150
rect 197400 74350 197600 74380
rect 197400 74150 197410 74350
rect 197480 74150 197520 74350
rect 197590 74150 197600 74350
rect 197400 74120 197600 74150
rect 197900 74350 198100 74380
rect 197900 74150 197910 74350
rect 197980 74150 198020 74350
rect 198090 74150 198100 74350
rect 197900 74120 198100 74150
rect 198400 74350 198600 74380
rect 198400 74150 198410 74350
rect 198480 74150 198520 74350
rect 198590 74150 198600 74350
rect 198400 74120 198600 74150
rect 198900 74350 199100 74380
rect 198900 74150 198910 74350
rect 198980 74150 199020 74350
rect 199090 74150 199100 74350
rect 198900 74120 199100 74150
rect 199400 74350 199600 74380
rect 199400 74150 199410 74350
rect 199480 74150 199520 74350
rect 199590 74150 199600 74350
rect 199400 74120 199600 74150
rect 199900 74350 200100 74380
rect 199900 74150 199910 74350
rect 199980 74150 200020 74350
rect 200090 74150 200100 74350
rect 199900 74120 200100 74150
rect 200400 74350 200600 74380
rect 200400 74150 200410 74350
rect 200480 74150 200520 74350
rect 200590 74150 200600 74350
rect 200400 74120 200600 74150
rect 200900 74350 201100 74380
rect 200900 74150 200910 74350
rect 200980 74150 201020 74350
rect 201090 74150 201100 74350
rect 200900 74120 201100 74150
rect 201400 74350 201600 74380
rect 201400 74150 201410 74350
rect 201480 74150 201520 74350
rect 201590 74150 201600 74350
rect 201400 74120 201600 74150
rect 201900 74350 202100 74380
rect 201900 74150 201910 74350
rect 201980 74150 202020 74350
rect 202090 74150 202100 74350
rect 201900 74120 202100 74150
rect 202400 74350 202600 74380
rect 202400 74150 202410 74350
rect 202480 74150 202520 74350
rect 202590 74150 202600 74350
rect 202400 74120 202600 74150
rect 202900 74350 203100 74380
rect 202900 74150 202910 74350
rect 202980 74150 203020 74350
rect 203090 74150 203100 74350
rect 202900 74120 203100 74150
rect 203400 74350 203600 74380
rect 203400 74150 203410 74350
rect 203480 74150 203520 74350
rect 203590 74150 203600 74350
rect 203400 74120 203600 74150
rect 203900 74350 204100 74380
rect 203900 74150 203910 74350
rect 203980 74150 204020 74350
rect 204090 74150 204100 74350
rect 203900 74120 204100 74150
rect 204400 74350 204600 74380
rect 204400 74150 204410 74350
rect 204480 74150 204520 74350
rect 204590 74150 204600 74350
rect 204400 74120 204600 74150
rect 204900 74350 205100 74380
rect 204900 74150 204910 74350
rect 204980 74150 205020 74350
rect 205090 74150 205100 74350
rect 204900 74120 205100 74150
rect 205400 74350 205600 74380
rect 205400 74150 205410 74350
rect 205480 74150 205520 74350
rect 205590 74150 205600 74350
rect 205400 74120 205600 74150
rect 205900 74350 206100 74380
rect 205900 74150 205910 74350
rect 205980 74150 206020 74350
rect 206090 74150 206100 74350
rect 205900 74120 206100 74150
rect 206400 74350 206600 74380
rect 206400 74150 206410 74350
rect 206480 74150 206520 74350
rect 206590 74150 206600 74350
rect 206400 74120 206600 74150
rect 206900 74350 207100 74380
rect 206900 74150 206910 74350
rect 206980 74150 207020 74350
rect 207090 74150 207100 74350
rect 206900 74120 207100 74150
rect 207400 74350 207600 74380
rect 207400 74150 207410 74350
rect 207480 74150 207520 74350
rect 207590 74150 207600 74350
rect 207400 74120 207600 74150
rect 207900 74350 208000 74380
rect 207900 74150 207910 74350
rect 207980 74150 208000 74350
rect 207900 74120 208000 74150
rect 196000 74100 196120 74120
rect 196380 74100 196620 74120
rect 196880 74100 197120 74120
rect 197380 74100 197620 74120
rect 197880 74100 198120 74120
rect 198380 74100 198620 74120
rect 198880 74100 199120 74120
rect 199380 74100 199620 74120
rect 199880 74100 200120 74120
rect 200380 74100 200620 74120
rect 200880 74100 201120 74120
rect 201380 74100 201620 74120
rect 201880 74100 202120 74120
rect 202380 74100 202620 74120
rect 202880 74100 203120 74120
rect 203380 74100 203620 74120
rect 203880 74100 204120 74120
rect 204380 74100 204620 74120
rect 204880 74100 205120 74120
rect 205380 74100 205620 74120
rect 205880 74100 206120 74120
rect 206380 74100 206620 74120
rect 206880 74100 207120 74120
rect 207380 74100 207620 74120
rect 207880 74100 208000 74120
rect 196000 74090 208000 74100
rect 196000 74020 196150 74090
rect 196350 74020 196650 74090
rect 196850 74020 197150 74090
rect 197350 74020 197650 74090
rect 197850 74020 198150 74090
rect 198350 74020 198650 74090
rect 198850 74020 199150 74090
rect 199350 74020 199650 74090
rect 199850 74020 200150 74090
rect 200350 74020 200650 74090
rect 200850 74020 201150 74090
rect 201350 74020 201650 74090
rect 201850 74020 202150 74090
rect 202350 74020 202650 74090
rect 202850 74020 203150 74090
rect 203350 74020 203650 74090
rect 203850 74020 204150 74090
rect 204350 74020 204650 74090
rect 204850 74020 205150 74090
rect 205350 74020 205650 74090
rect 205850 74020 206150 74090
rect 206350 74020 206650 74090
rect 206850 74020 207150 74090
rect 207350 74020 207650 74090
rect 207850 74020 208000 74090
rect 196000 73980 208000 74020
rect 196000 73910 196150 73980
rect 196350 73910 196650 73980
rect 196850 73910 197150 73980
rect 197350 73910 197650 73980
rect 197850 73910 198150 73980
rect 198350 73910 198650 73980
rect 198850 73910 199150 73980
rect 199350 73910 199650 73980
rect 199850 73910 200150 73980
rect 200350 73910 200650 73980
rect 200850 73910 201150 73980
rect 201350 73910 201650 73980
rect 201850 73910 202150 73980
rect 202350 73910 202650 73980
rect 202850 73910 203150 73980
rect 203350 73910 203650 73980
rect 203850 73910 204150 73980
rect 204350 73910 204650 73980
rect 204850 73910 205150 73980
rect 205350 73910 205650 73980
rect 205850 73910 206150 73980
rect 206350 73910 206650 73980
rect 206850 73910 207150 73980
rect 207350 73910 207650 73980
rect 207850 73910 208000 73980
rect 196000 73900 208000 73910
rect 196000 73880 196120 73900
rect 196380 73880 196620 73900
rect 196880 73880 197120 73900
rect 197380 73880 197620 73900
rect 197880 73880 198120 73900
rect 198380 73880 198620 73900
rect 198880 73880 199120 73900
rect 199380 73880 199620 73900
rect 199880 73880 200120 73900
rect 200380 73880 200620 73900
rect 200880 73880 201120 73900
rect 201380 73880 201620 73900
rect 201880 73880 202120 73900
rect 202380 73880 202620 73900
rect 202880 73880 203120 73900
rect 203380 73880 203620 73900
rect 203880 73880 204120 73900
rect 204380 73880 204620 73900
rect 204880 73880 205120 73900
rect 205380 73880 205620 73900
rect 205880 73880 206120 73900
rect 206380 73880 206620 73900
rect 206880 73880 207120 73900
rect 207380 73880 207620 73900
rect 207880 73880 208000 73900
rect 196000 73850 196100 73880
rect 196000 73650 196020 73850
rect 196090 73650 196100 73850
rect 196000 73620 196100 73650
rect 196400 73850 196600 73880
rect 196400 73650 196410 73850
rect 196480 73650 196520 73850
rect 196590 73650 196600 73850
rect 196400 73620 196600 73650
rect 196900 73850 197100 73880
rect 196900 73650 196910 73850
rect 196980 73650 197020 73850
rect 197090 73650 197100 73850
rect 196900 73620 197100 73650
rect 197400 73850 197600 73880
rect 197400 73650 197410 73850
rect 197480 73650 197520 73850
rect 197590 73650 197600 73850
rect 197400 73620 197600 73650
rect 197900 73850 198100 73880
rect 197900 73650 197910 73850
rect 197980 73650 198020 73850
rect 198090 73650 198100 73850
rect 197900 73620 198100 73650
rect 198400 73850 198600 73880
rect 198400 73650 198410 73850
rect 198480 73650 198520 73850
rect 198590 73650 198600 73850
rect 198400 73620 198600 73650
rect 198900 73850 199100 73880
rect 198900 73650 198910 73850
rect 198980 73650 199020 73850
rect 199090 73650 199100 73850
rect 198900 73620 199100 73650
rect 199400 73850 199600 73880
rect 199400 73650 199410 73850
rect 199480 73650 199520 73850
rect 199590 73650 199600 73850
rect 199400 73620 199600 73650
rect 199900 73850 200100 73880
rect 199900 73650 199910 73850
rect 199980 73650 200020 73850
rect 200090 73650 200100 73850
rect 199900 73620 200100 73650
rect 200400 73850 200600 73880
rect 200400 73650 200410 73850
rect 200480 73650 200520 73850
rect 200590 73650 200600 73850
rect 200400 73620 200600 73650
rect 200900 73850 201100 73880
rect 200900 73650 200910 73850
rect 200980 73650 201020 73850
rect 201090 73650 201100 73850
rect 200900 73620 201100 73650
rect 201400 73850 201600 73880
rect 201400 73650 201410 73850
rect 201480 73650 201520 73850
rect 201590 73650 201600 73850
rect 201400 73620 201600 73650
rect 201900 73850 202100 73880
rect 201900 73650 201910 73850
rect 201980 73650 202020 73850
rect 202090 73650 202100 73850
rect 201900 73620 202100 73650
rect 202400 73850 202600 73880
rect 202400 73650 202410 73850
rect 202480 73650 202520 73850
rect 202590 73650 202600 73850
rect 202400 73620 202600 73650
rect 202900 73850 203100 73880
rect 202900 73650 202910 73850
rect 202980 73650 203020 73850
rect 203090 73650 203100 73850
rect 202900 73620 203100 73650
rect 203400 73850 203600 73880
rect 203400 73650 203410 73850
rect 203480 73650 203520 73850
rect 203590 73650 203600 73850
rect 203400 73620 203600 73650
rect 203900 73850 204100 73880
rect 203900 73650 203910 73850
rect 203980 73650 204020 73850
rect 204090 73650 204100 73850
rect 203900 73620 204100 73650
rect 204400 73850 204600 73880
rect 204400 73650 204410 73850
rect 204480 73650 204520 73850
rect 204590 73650 204600 73850
rect 204400 73620 204600 73650
rect 204900 73850 205100 73880
rect 204900 73650 204910 73850
rect 204980 73650 205020 73850
rect 205090 73650 205100 73850
rect 204900 73620 205100 73650
rect 205400 73850 205600 73880
rect 205400 73650 205410 73850
rect 205480 73650 205520 73850
rect 205590 73650 205600 73850
rect 205400 73620 205600 73650
rect 205900 73850 206100 73880
rect 205900 73650 205910 73850
rect 205980 73650 206020 73850
rect 206090 73650 206100 73850
rect 205900 73620 206100 73650
rect 206400 73850 206600 73880
rect 206400 73650 206410 73850
rect 206480 73650 206520 73850
rect 206590 73650 206600 73850
rect 206400 73620 206600 73650
rect 206900 73850 207100 73880
rect 206900 73650 206910 73850
rect 206980 73650 207020 73850
rect 207090 73650 207100 73850
rect 206900 73620 207100 73650
rect 207400 73850 207600 73880
rect 207400 73650 207410 73850
rect 207480 73650 207520 73850
rect 207590 73650 207600 73850
rect 207400 73620 207600 73650
rect 207900 73850 208000 73880
rect 207900 73650 207910 73850
rect 207980 73650 208000 73850
rect 207900 73620 208000 73650
rect 196000 73600 196120 73620
rect 196380 73600 196620 73620
rect 196880 73600 197120 73620
rect 197380 73600 197620 73620
rect 197880 73600 198120 73620
rect 198380 73600 198620 73620
rect 198880 73600 199120 73620
rect 199380 73600 199620 73620
rect 199880 73600 200120 73620
rect 200380 73600 200620 73620
rect 200880 73600 201120 73620
rect 201380 73600 201620 73620
rect 201880 73600 202120 73620
rect 202380 73600 202620 73620
rect 202880 73600 203120 73620
rect 203380 73600 203620 73620
rect 203880 73600 204120 73620
rect 204380 73600 204620 73620
rect 204880 73600 205120 73620
rect 205380 73600 205620 73620
rect 205880 73600 206120 73620
rect 206380 73600 206620 73620
rect 206880 73600 207120 73620
rect 207380 73600 207620 73620
rect 207880 73600 208000 73620
rect 196000 73590 208000 73600
rect 196000 73520 196150 73590
rect 196350 73520 196650 73590
rect 196850 73520 197150 73590
rect 197350 73520 197650 73590
rect 197850 73520 198150 73590
rect 198350 73520 198650 73590
rect 198850 73520 199150 73590
rect 199350 73520 199650 73590
rect 199850 73520 200150 73590
rect 200350 73520 200650 73590
rect 200850 73520 201150 73590
rect 201350 73520 201650 73590
rect 201850 73520 202150 73590
rect 202350 73520 202650 73590
rect 202850 73520 203150 73590
rect 203350 73520 203650 73590
rect 203850 73520 204150 73590
rect 204350 73520 204650 73590
rect 204850 73520 205150 73590
rect 205350 73520 205650 73590
rect 205850 73520 206150 73590
rect 206350 73520 206650 73590
rect 206850 73520 207150 73590
rect 207350 73520 207650 73590
rect 207850 73520 208000 73590
rect 196000 73480 208000 73520
rect 196000 73410 196150 73480
rect 196350 73410 196650 73480
rect 196850 73410 197150 73480
rect 197350 73410 197650 73480
rect 197850 73410 198150 73480
rect 198350 73410 198650 73480
rect 198850 73410 199150 73480
rect 199350 73410 199650 73480
rect 199850 73410 200150 73480
rect 200350 73410 200650 73480
rect 200850 73410 201150 73480
rect 201350 73410 201650 73480
rect 201850 73410 202150 73480
rect 202350 73410 202650 73480
rect 202850 73410 203150 73480
rect 203350 73410 203650 73480
rect 203850 73410 204150 73480
rect 204350 73410 204650 73480
rect 204850 73410 205150 73480
rect 205350 73410 205650 73480
rect 205850 73410 206150 73480
rect 206350 73410 206650 73480
rect 206850 73410 207150 73480
rect 207350 73410 207650 73480
rect 207850 73410 208000 73480
rect 196000 73400 208000 73410
rect 196000 73380 196120 73400
rect 196380 73380 196620 73400
rect 196880 73380 197120 73400
rect 197380 73380 197620 73400
rect 197880 73380 198120 73400
rect 198380 73380 198620 73400
rect 198880 73380 199120 73400
rect 199380 73380 199620 73400
rect 199880 73380 200120 73400
rect 200380 73380 200620 73400
rect 200880 73380 201120 73400
rect 201380 73380 201620 73400
rect 201880 73380 202120 73400
rect 202380 73380 202620 73400
rect 202880 73380 203120 73400
rect 203380 73380 203620 73400
rect 203880 73380 204120 73400
rect 204380 73380 204620 73400
rect 204880 73380 205120 73400
rect 205380 73380 205620 73400
rect 205880 73380 206120 73400
rect 206380 73380 206620 73400
rect 206880 73380 207120 73400
rect 207380 73380 207620 73400
rect 207880 73380 208000 73400
rect 196000 73350 196100 73380
rect 196000 73150 196020 73350
rect 196090 73150 196100 73350
rect 196000 73120 196100 73150
rect 196400 73350 196600 73380
rect 196400 73150 196410 73350
rect 196480 73150 196520 73350
rect 196590 73150 196600 73350
rect 196400 73120 196600 73150
rect 196900 73350 197100 73380
rect 196900 73150 196910 73350
rect 196980 73150 197020 73350
rect 197090 73150 197100 73350
rect 196900 73120 197100 73150
rect 197400 73350 197600 73380
rect 197400 73150 197410 73350
rect 197480 73150 197520 73350
rect 197590 73150 197600 73350
rect 197400 73120 197600 73150
rect 197900 73350 198100 73380
rect 197900 73150 197910 73350
rect 197980 73150 198020 73350
rect 198090 73150 198100 73350
rect 197900 73120 198100 73150
rect 198400 73350 198600 73380
rect 198400 73150 198410 73350
rect 198480 73150 198520 73350
rect 198590 73150 198600 73350
rect 198400 73120 198600 73150
rect 198900 73350 199100 73380
rect 198900 73150 198910 73350
rect 198980 73150 199020 73350
rect 199090 73150 199100 73350
rect 198900 73120 199100 73150
rect 199400 73350 199600 73380
rect 199400 73150 199410 73350
rect 199480 73150 199520 73350
rect 199590 73150 199600 73350
rect 199400 73120 199600 73150
rect 199900 73350 200100 73380
rect 199900 73150 199910 73350
rect 199980 73150 200020 73350
rect 200090 73150 200100 73350
rect 199900 73120 200100 73150
rect 200400 73350 200600 73380
rect 200400 73150 200410 73350
rect 200480 73150 200520 73350
rect 200590 73150 200600 73350
rect 200400 73120 200600 73150
rect 200900 73350 201100 73380
rect 200900 73150 200910 73350
rect 200980 73150 201020 73350
rect 201090 73150 201100 73350
rect 200900 73120 201100 73150
rect 201400 73350 201600 73380
rect 201400 73150 201410 73350
rect 201480 73150 201520 73350
rect 201590 73150 201600 73350
rect 201400 73120 201600 73150
rect 201900 73350 202100 73380
rect 201900 73150 201910 73350
rect 201980 73150 202020 73350
rect 202090 73150 202100 73350
rect 201900 73120 202100 73150
rect 202400 73350 202600 73380
rect 202400 73150 202410 73350
rect 202480 73150 202520 73350
rect 202590 73150 202600 73350
rect 202400 73120 202600 73150
rect 202900 73350 203100 73380
rect 202900 73150 202910 73350
rect 202980 73150 203020 73350
rect 203090 73150 203100 73350
rect 202900 73120 203100 73150
rect 203400 73350 203600 73380
rect 203400 73150 203410 73350
rect 203480 73150 203520 73350
rect 203590 73150 203600 73350
rect 203400 73120 203600 73150
rect 203900 73350 204100 73380
rect 203900 73150 203910 73350
rect 203980 73150 204020 73350
rect 204090 73150 204100 73350
rect 203900 73120 204100 73150
rect 204400 73350 204600 73380
rect 204400 73150 204410 73350
rect 204480 73150 204520 73350
rect 204590 73150 204600 73350
rect 204400 73120 204600 73150
rect 204900 73350 205100 73380
rect 204900 73150 204910 73350
rect 204980 73150 205020 73350
rect 205090 73150 205100 73350
rect 204900 73120 205100 73150
rect 205400 73350 205600 73380
rect 205400 73150 205410 73350
rect 205480 73150 205520 73350
rect 205590 73150 205600 73350
rect 205400 73120 205600 73150
rect 205900 73350 206100 73380
rect 205900 73150 205910 73350
rect 205980 73150 206020 73350
rect 206090 73150 206100 73350
rect 205900 73120 206100 73150
rect 206400 73350 206600 73380
rect 206400 73150 206410 73350
rect 206480 73150 206520 73350
rect 206590 73150 206600 73350
rect 206400 73120 206600 73150
rect 206900 73350 207100 73380
rect 206900 73150 206910 73350
rect 206980 73150 207020 73350
rect 207090 73150 207100 73350
rect 206900 73120 207100 73150
rect 207400 73350 207600 73380
rect 207400 73150 207410 73350
rect 207480 73150 207520 73350
rect 207590 73150 207600 73350
rect 207400 73120 207600 73150
rect 207900 73350 208000 73380
rect 207900 73150 207910 73350
rect 207980 73150 208000 73350
rect 207900 73120 208000 73150
rect 196000 73100 196120 73120
rect 196380 73100 196620 73120
rect 196880 73100 197120 73120
rect 197380 73100 197620 73120
rect 197880 73100 198120 73120
rect 198380 73100 198620 73120
rect 198880 73100 199120 73120
rect 199380 73100 199620 73120
rect 199880 73100 200120 73120
rect 200380 73100 200620 73120
rect 200880 73100 201120 73120
rect 201380 73100 201620 73120
rect 201880 73100 202120 73120
rect 202380 73100 202620 73120
rect 202880 73100 203120 73120
rect 203380 73100 203620 73120
rect 203880 73100 204120 73120
rect 204380 73100 204620 73120
rect 204880 73100 205120 73120
rect 205380 73100 205620 73120
rect 205880 73100 206120 73120
rect 206380 73100 206620 73120
rect 206880 73100 207120 73120
rect 207380 73100 207620 73120
rect 207880 73100 208000 73120
rect 196000 73090 208000 73100
rect 196000 73020 196150 73090
rect 196350 73020 196650 73090
rect 196850 73020 197150 73090
rect 197350 73020 197650 73090
rect 197850 73020 198150 73090
rect 198350 73020 198650 73090
rect 198850 73020 199150 73090
rect 199350 73020 199650 73090
rect 199850 73020 200150 73090
rect 200350 73020 200650 73090
rect 200850 73020 201150 73090
rect 201350 73020 201650 73090
rect 201850 73020 202150 73090
rect 202350 73020 202650 73090
rect 202850 73020 203150 73090
rect 203350 73020 203650 73090
rect 203850 73020 204150 73090
rect 204350 73020 204650 73090
rect 204850 73020 205150 73090
rect 205350 73020 205650 73090
rect 205850 73020 206150 73090
rect 206350 73020 206650 73090
rect 206850 73020 207150 73090
rect 207350 73020 207650 73090
rect 207850 73020 208000 73090
rect 196000 72980 208000 73020
rect 196000 72910 196150 72980
rect 196350 72910 196650 72980
rect 196850 72910 197150 72980
rect 197350 72910 197650 72980
rect 197850 72910 198150 72980
rect 198350 72910 198650 72980
rect 198850 72910 199150 72980
rect 199350 72910 199650 72980
rect 199850 72910 200150 72980
rect 200350 72910 200650 72980
rect 200850 72910 201150 72980
rect 201350 72910 201650 72980
rect 201850 72910 202150 72980
rect 202350 72910 202650 72980
rect 202850 72910 203150 72980
rect 203350 72910 203650 72980
rect 203850 72910 204150 72980
rect 204350 72910 204650 72980
rect 204850 72910 205150 72980
rect 205350 72910 205650 72980
rect 205850 72910 206150 72980
rect 206350 72910 206650 72980
rect 206850 72910 207150 72980
rect 207350 72910 207650 72980
rect 207850 72910 208000 72980
rect 196000 72900 208000 72910
rect 196000 72880 196120 72900
rect 196380 72880 196620 72900
rect 196880 72880 197120 72900
rect 197380 72880 197620 72900
rect 197880 72880 198120 72900
rect 198380 72880 198620 72900
rect 198880 72880 199120 72900
rect 199380 72880 199620 72900
rect 199880 72880 200120 72900
rect 200380 72880 200620 72900
rect 200880 72880 201120 72900
rect 201380 72880 201620 72900
rect 201880 72880 202120 72900
rect 202380 72880 202620 72900
rect 202880 72880 203120 72900
rect 203380 72880 203620 72900
rect 203880 72880 204120 72900
rect 204380 72880 204620 72900
rect 204880 72880 205120 72900
rect 205380 72880 205620 72900
rect 205880 72880 206120 72900
rect 206380 72880 206620 72900
rect 206880 72880 207120 72900
rect 207380 72880 207620 72900
rect 207880 72880 208000 72900
rect 196000 72850 196100 72880
rect 196000 72650 196020 72850
rect 196090 72650 196100 72850
rect 196000 72620 196100 72650
rect 196400 72850 196600 72880
rect 196400 72650 196410 72850
rect 196480 72650 196520 72850
rect 196590 72650 196600 72850
rect 196400 72620 196600 72650
rect 196900 72850 197100 72880
rect 196900 72650 196910 72850
rect 196980 72650 197020 72850
rect 197090 72650 197100 72850
rect 196900 72620 197100 72650
rect 197400 72850 197600 72880
rect 197400 72650 197410 72850
rect 197480 72650 197520 72850
rect 197590 72650 197600 72850
rect 197400 72620 197600 72650
rect 197900 72850 198100 72880
rect 197900 72650 197910 72850
rect 197980 72650 198020 72850
rect 198090 72650 198100 72850
rect 197900 72620 198100 72650
rect 198400 72850 198600 72880
rect 198400 72650 198410 72850
rect 198480 72650 198520 72850
rect 198590 72650 198600 72850
rect 198400 72620 198600 72650
rect 198900 72850 199100 72880
rect 198900 72650 198910 72850
rect 198980 72650 199020 72850
rect 199090 72650 199100 72850
rect 198900 72620 199100 72650
rect 199400 72850 199600 72880
rect 199400 72650 199410 72850
rect 199480 72650 199520 72850
rect 199590 72650 199600 72850
rect 199400 72620 199600 72650
rect 199900 72850 200100 72880
rect 199900 72650 199910 72850
rect 199980 72650 200020 72850
rect 200090 72650 200100 72850
rect 199900 72620 200100 72650
rect 200400 72850 200600 72880
rect 200400 72650 200410 72850
rect 200480 72650 200520 72850
rect 200590 72650 200600 72850
rect 200400 72620 200600 72650
rect 200900 72850 201100 72880
rect 200900 72650 200910 72850
rect 200980 72650 201020 72850
rect 201090 72650 201100 72850
rect 200900 72620 201100 72650
rect 201400 72850 201600 72880
rect 201400 72650 201410 72850
rect 201480 72650 201520 72850
rect 201590 72650 201600 72850
rect 201400 72620 201600 72650
rect 201900 72850 202100 72880
rect 201900 72650 201910 72850
rect 201980 72650 202020 72850
rect 202090 72650 202100 72850
rect 201900 72620 202100 72650
rect 202400 72850 202600 72880
rect 202400 72650 202410 72850
rect 202480 72650 202520 72850
rect 202590 72650 202600 72850
rect 202400 72620 202600 72650
rect 202900 72850 203100 72880
rect 202900 72650 202910 72850
rect 202980 72650 203020 72850
rect 203090 72650 203100 72850
rect 202900 72620 203100 72650
rect 203400 72850 203600 72880
rect 203400 72650 203410 72850
rect 203480 72650 203520 72850
rect 203590 72650 203600 72850
rect 203400 72620 203600 72650
rect 203900 72850 204100 72880
rect 203900 72650 203910 72850
rect 203980 72650 204020 72850
rect 204090 72650 204100 72850
rect 203900 72620 204100 72650
rect 204400 72850 204600 72880
rect 204400 72650 204410 72850
rect 204480 72650 204520 72850
rect 204590 72650 204600 72850
rect 204400 72620 204600 72650
rect 204900 72850 205100 72880
rect 204900 72650 204910 72850
rect 204980 72650 205020 72850
rect 205090 72650 205100 72850
rect 204900 72620 205100 72650
rect 205400 72850 205600 72880
rect 205400 72650 205410 72850
rect 205480 72650 205520 72850
rect 205590 72650 205600 72850
rect 205400 72620 205600 72650
rect 205900 72850 206100 72880
rect 205900 72650 205910 72850
rect 205980 72650 206020 72850
rect 206090 72650 206100 72850
rect 205900 72620 206100 72650
rect 206400 72850 206600 72880
rect 206400 72650 206410 72850
rect 206480 72650 206520 72850
rect 206590 72650 206600 72850
rect 206400 72620 206600 72650
rect 206900 72850 207100 72880
rect 206900 72650 206910 72850
rect 206980 72650 207020 72850
rect 207090 72650 207100 72850
rect 206900 72620 207100 72650
rect 207400 72850 207600 72880
rect 207400 72650 207410 72850
rect 207480 72650 207520 72850
rect 207590 72650 207600 72850
rect 207400 72620 207600 72650
rect 207900 72850 208000 72880
rect 207900 72650 207910 72850
rect 207980 72650 208000 72850
rect 207900 72620 208000 72650
rect 196000 72600 196120 72620
rect 196380 72600 196620 72620
rect 196880 72600 197120 72620
rect 197380 72600 197620 72620
rect 197880 72600 198120 72620
rect 198380 72600 198620 72620
rect 198880 72600 199120 72620
rect 199380 72600 199620 72620
rect 199880 72600 200120 72620
rect 200380 72600 200620 72620
rect 200880 72600 201120 72620
rect 201380 72600 201620 72620
rect 201880 72600 202120 72620
rect 202380 72600 202620 72620
rect 202880 72600 203120 72620
rect 203380 72600 203620 72620
rect 203880 72600 204120 72620
rect 204380 72600 204620 72620
rect 204880 72600 205120 72620
rect 205380 72600 205620 72620
rect 205880 72600 206120 72620
rect 206380 72600 206620 72620
rect 206880 72600 207120 72620
rect 207380 72600 207620 72620
rect 207880 72600 208000 72620
rect 196000 72590 208000 72600
rect 196000 72520 196150 72590
rect 196350 72520 196650 72590
rect 196850 72520 197150 72590
rect 197350 72520 197650 72590
rect 197850 72520 198150 72590
rect 198350 72520 198650 72590
rect 198850 72520 199150 72590
rect 199350 72520 199650 72590
rect 199850 72520 200150 72590
rect 200350 72520 200650 72590
rect 200850 72520 201150 72590
rect 201350 72520 201650 72590
rect 201850 72520 202150 72590
rect 202350 72520 202650 72590
rect 202850 72520 203150 72590
rect 203350 72520 203650 72590
rect 203850 72520 204150 72590
rect 204350 72520 204650 72590
rect 204850 72520 205150 72590
rect 205350 72520 205650 72590
rect 205850 72520 206150 72590
rect 206350 72520 206650 72590
rect 206850 72520 207150 72590
rect 207350 72520 207650 72590
rect 207850 72520 208000 72590
rect 196000 72480 208000 72520
rect 196000 72410 196150 72480
rect 196350 72410 196650 72480
rect 196850 72410 197150 72480
rect 197350 72410 197650 72480
rect 197850 72410 198150 72480
rect 198350 72410 198650 72480
rect 198850 72410 199150 72480
rect 199350 72410 199650 72480
rect 199850 72410 200150 72480
rect 200350 72410 200650 72480
rect 200850 72410 201150 72480
rect 201350 72410 201650 72480
rect 201850 72410 202150 72480
rect 202350 72410 202650 72480
rect 202850 72410 203150 72480
rect 203350 72410 203650 72480
rect 203850 72410 204150 72480
rect 204350 72410 204650 72480
rect 204850 72410 205150 72480
rect 205350 72410 205650 72480
rect 205850 72410 206150 72480
rect 206350 72410 206650 72480
rect 206850 72410 207150 72480
rect 207350 72410 207650 72480
rect 207850 72410 208000 72480
rect 196000 72400 208000 72410
rect 196000 72380 196120 72400
rect 196380 72380 196620 72400
rect 196880 72380 197120 72400
rect 197380 72380 197620 72400
rect 197880 72380 198120 72400
rect 198380 72380 198620 72400
rect 198880 72380 199120 72400
rect 199380 72380 199620 72400
rect 199880 72380 200120 72400
rect 200380 72380 200620 72400
rect 200880 72380 201120 72400
rect 201380 72380 201620 72400
rect 201880 72380 202120 72400
rect 202380 72380 202620 72400
rect 202880 72380 203120 72400
rect 203380 72380 203620 72400
rect 203880 72380 204120 72400
rect 204380 72380 204620 72400
rect 204880 72380 205120 72400
rect 205380 72380 205620 72400
rect 205880 72380 206120 72400
rect 206380 72380 206620 72400
rect 206880 72380 207120 72400
rect 207380 72380 207620 72400
rect 207880 72380 208000 72400
rect 196000 72350 196100 72380
rect 196000 72150 196020 72350
rect 196090 72150 196100 72350
rect 196000 72120 196100 72150
rect 196400 72350 196600 72380
rect 196400 72150 196410 72350
rect 196480 72150 196520 72350
rect 196590 72150 196600 72350
rect 196400 72120 196600 72150
rect 196900 72350 197100 72380
rect 196900 72150 196910 72350
rect 196980 72150 197020 72350
rect 197090 72150 197100 72350
rect 196900 72120 197100 72150
rect 197400 72350 197600 72380
rect 197400 72150 197410 72350
rect 197480 72150 197520 72350
rect 197590 72150 197600 72350
rect 197400 72120 197600 72150
rect 197900 72350 198100 72380
rect 197900 72150 197910 72350
rect 197980 72150 198020 72350
rect 198090 72150 198100 72350
rect 197900 72120 198100 72150
rect 198400 72350 198600 72380
rect 198400 72150 198410 72350
rect 198480 72150 198520 72350
rect 198590 72150 198600 72350
rect 198400 72120 198600 72150
rect 198900 72350 199100 72380
rect 198900 72150 198910 72350
rect 198980 72150 199020 72350
rect 199090 72150 199100 72350
rect 198900 72120 199100 72150
rect 199400 72350 199600 72380
rect 199400 72150 199410 72350
rect 199480 72150 199520 72350
rect 199590 72150 199600 72350
rect 199400 72120 199600 72150
rect 199900 72350 200100 72380
rect 199900 72150 199910 72350
rect 199980 72150 200020 72350
rect 200090 72150 200100 72350
rect 199900 72120 200100 72150
rect 200400 72350 200600 72380
rect 200400 72150 200410 72350
rect 200480 72150 200520 72350
rect 200590 72150 200600 72350
rect 200400 72120 200600 72150
rect 200900 72350 201100 72380
rect 200900 72150 200910 72350
rect 200980 72150 201020 72350
rect 201090 72150 201100 72350
rect 200900 72120 201100 72150
rect 201400 72350 201600 72380
rect 201400 72150 201410 72350
rect 201480 72150 201520 72350
rect 201590 72150 201600 72350
rect 201400 72120 201600 72150
rect 201900 72350 202100 72380
rect 201900 72150 201910 72350
rect 201980 72150 202020 72350
rect 202090 72150 202100 72350
rect 201900 72120 202100 72150
rect 202400 72350 202600 72380
rect 202400 72150 202410 72350
rect 202480 72150 202520 72350
rect 202590 72150 202600 72350
rect 202400 72120 202600 72150
rect 202900 72350 203100 72380
rect 202900 72150 202910 72350
rect 202980 72150 203020 72350
rect 203090 72150 203100 72350
rect 202900 72120 203100 72150
rect 203400 72350 203600 72380
rect 203400 72150 203410 72350
rect 203480 72150 203520 72350
rect 203590 72150 203600 72350
rect 203400 72120 203600 72150
rect 203900 72350 204100 72380
rect 203900 72150 203910 72350
rect 203980 72150 204020 72350
rect 204090 72150 204100 72350
rect 203900 72120 204100 72150
rect 204400 72350 204600 72380
rect 204400 72150 204410 72350
rect 204480 72150 204520 72350
rect 204590 72150 204600 72350
rect 204400 72120 204600 72150
rect 204900 72350 205100 72380
rect 204900 72150 204910 72350
rect 204980 72150 205020 72350
rect 205090 72150 205100 72350
rect 204900 72120 205100 72150
rect 205400 72350 205600 72380
rect 205400 72150 205410 72350
rect 205480 72150 205520 72350
rect 205590 72150 205600 72350
rect 205400 72120 205600 72150
rect 205900 72350 206100 72380
rect 205900 72150 205910 72350
rect 205980 72150 206020 72350
rect 206090 72150 206100 72350
rect 205900 72120 206100 72150
rect 206400 72350 206600 72380
rect 206400 72150 206410 72350
rect 206480 72150 206520 72350
rect 206590 72150 206600 72350
rect 206400 72120 206600 72150
rect 206900 72350 207100 72380
rect 206900 72150 206910 72350
rect 206980 72150 207020 72350
rect 207090 72150 207100 72350
rect 206900 72120 207100 72150
rect 207400 72350 207600 72380
rect 207400 72150 207410 72350
rect 207480 72150 207520 72350
rect 207590 72150 207600 72350
rect 207400 72120 207600 72150
rect 207900 72350 208000 72380
rect 207900 72150 207910 72350
rect 207980 72150 208000 72350
rect 207900 72120 208000 72150
rect 196000 72100 196120 72120
rect 196380 72100 196620 72120
rect 196880 72100 197120 72120
rect 197380 72100 197620 72120
rect 197880 72100 198120 72120
rect 198380 72100 198620 72120
rect 198880 72100 199120 72120
rect 199380 72100 199620 72120
rect 199880 72100 200120 72120
rect 200380 72100 200620 72120
rect 200880 72100 201120 72120
rect 201380 72100 201620 72120
rect 201880 72100 202120 72120
rect 202380 72100 202620 72120
rect 202880 72100 203120 72120
rect 203380 72100 203620 72120
rect 203880 72100 204120 72120
rect 204380 72100 204620 72120
rect 204880 72100 205120 72120
rect 205380 72100 205620 72120
rect 205880 72100 206120 72120
rect 206380 72100 206620 72120
rect 206880 72100 207120 72120
rect 207380 72100 207620 72120
rect 207880 72100 208000 72120
rect 196000 72090 208000 72100
rect 196000 72020 196150 72090
rect 196350 72020 196650 72090
rect 196850 72020 197150 72090
rect 197350 72020 197650 72090
rect 197850 72020 198150 72090
rect 198350 72020 198650 72090
rect 198850 72020 199150 72090
rect 199350 72020 199650 72090
rect 199850 72020 200150 72090
rect 200350 72020 200650 72090
rect 200850 72020 201150 72090
rect 201350 72020 201650 72090
rect 201850 72020 202150 72090
rect 202350 72020 202650 72090
rect 202850 72020 203150 72090
rect 203350 72020 203650 72090
rect 203850 72020 204150 72090
rect 204350 72020 204650 72090
rect 204850 72020 205150 72090
rect 205350 72020 205650 72090
rect 205850 72020 206150 72090
rect 206350 72020 206650 72090
rect 206850 72020 207150 72090
rect 207350 72020 207650 72090
rect 207850 72020 208000 72090
rect 196000 71980 208000 72020
rect 196000 71910 196150 71980
rect 196350 71910 196650 71980
rect 196850 71910 197150 71980
rect 197350 71910 197650 71980
rect 197850 71910 198150 71980
rect 198350 71910 198650 71980
rect 198850 71910 199150 71980
rect 199350 71910 199650 71980
rect 199850 71910 200150 71980
rect 200350 71910 200650 71980
rect 200850 71910 201150 71980
rect 201350 71910 201650 71980
rect 201850 71910 202150 71980
rect 202350 71910 202650 71980
rect 202850 71910 203150 71980
rect 203350 71910 203650 71980
rect 203850 71910 204150 71980
rect 204350 71910 204650 71980
rect 204850 71910 205150 71980
rect 205350 71910 205650 71980
rect 205850 71910 206150 71980
rect 206350 71910 206650 71980
rect 206850 71910 207150 71980
rect 207350 71910 207650 71980
rect 207850 71910 208000 71980
rect 196000 71900 208000 71910
rect 196000 71880 196120 71900
rect 196380 71880 196620 71900
rect 196880 71880 197120 71900
rect 197380 71880 197620 71900
rect 197880 71880 198120 71900
rect 198380 71880 198620 71900
rect 198880 71880 199120 71900
rect 199380 71880 199620 71900
rect 199880 71880 200120 71900
rect 200380 71880 200620 71900
rect 200880 71880 201120 71900
rect 201380 71880 201620 71900
rect 201880 71880 202120 71900
rect 202380 71880 202620 71900
rect 202880 71880 203120 71900
rect 203380 71880 203620 71900
rect 203880 71880 204120 71900
rect 204380 71880 204620 71900
rect 204880 71880 205120 71900
rect 205380 71880 205620 71900
rect 205880 71880 206120 71900
rect 206380 71880 206620 71900
rect 206880 71880 207120 71900
rect 207380 71880 207620 71900
rect 207880 71880 208000 71900
rect 196000 71850 196100 71880
rect 196000 71650 196020 71850
rect 196090 71650 196100 71850
rect 196000 71620 196100 71650
rect 196400 71850 196600 71880
rect 196400 71650 196410 71850
rect 196480 71650 196520 71850
rect 196590 71650 196600 71850
rect 196400 71620 196600 71650
rect 196900 71850 197100 71880
rect 196900 71650 196910 71850
rect 196980 71650 197020 71850
rect 197090 71650 197100 71850
rect 196900 71620 197100 71650
rect 197400 71850 197600 71880
rect 197400 71650 197410 71850
rect 197480 71650 197520 71850
rect 197590 71650 197600 71850
rect 197400 71620 197600 71650
rect 197900 71850 198100 71880
rect 197900 71650 197910 71850
rect 197980 71650 198020 71850
rect 198090 71650 198100 71850
rect 197900 71620 198100 71650
rect 198400 71850 198600 71880
rect 198400 71650 198410 71850
rect 198480 71650 198520 71850
rect 198590 71650 198600 71850
rect 198400 71620 198600 71650
rect 198900 71850 199100 71880
rect 198900 71650 198910 71850
rect 198980 71650 199020 71850
rect 199090 71650 199100 71850
rect 198900 71620 199100 71650
rect 199400 71850 199600 71880
rect 199400 71650 199410 71850
rect 199480 71650 199520 71850
rect 199590 71650 199600 71850
rect 199400 71620 199600 71650
rect 199900 71850 200100 71880
rect 199900 71650 199910 71850
rect 199980 71650 200020 71850
rect 200090 71650 200100 71850
rect 199900 71620 200100 71650
rect 200400 71850 200600 71880
rect 200400 71650 200410 71850
rect 200480 71650 200520 71850
rect 200590 71650 200600 71850
rect 200400 71620 200600 71650
rect 200900 71850 201100 71880
rect 200900 71650 200910 71850
rect 200980 71650 201020 71850
rect 201090 71650 201100 71850
rect 200900 71620 201100 71650
rect 201400 71850 201600 71880
rect 201400 71650 201410 71850
rect 201480 71650 201520 71850
rect 201590 71650 201600 71850
rect 201400 71620 201600 71650
rect 201900 71850 202100 71880
rect 201900 71650 201910 71850
rect 201980 71650 202020 71850
rect 202090 71650 202100 71850
rect 201900 71620 202100 71650
rect 202400 71850 202600 71880
rect 202400 71650 202410 71850
rect 202480 71650 202520 71850
rect 202590 71650 202600 71850
rect 202400 71620 202600 71650
rect 202900 71850 203100 71880
rect 202900 71650 202910 71850
rect 202980 71650 203020 71850
rect 203090 71650 203100 71850
rect 202900 71620 203100 71650
rect 203400 71850 203600 71880
rect 203400 71650 203410 71850
rect 203480 71650 203520 71850
rect 203590 71650 203600 71850
rect 203400 71620 203600 71650
rect 203900 71850 204100 71880
rect 203900 71650 203910 71850
rect 203980 71650 204020 71850
rect 204090 71650 204100 71850
rect 203900 71620 204100 71650
rect 204400 71850 204600 71880
rect 204400 71650 204410 71850
rect 204480 71650 204520 71850
rect 204590 71650 204600 71850
rect 204400 71620 204600 71650
rect 204900 71850 205100 71880
rect 204900 71650 204910 71850
rect 204980 71650 205020 71850
rect 205090 71650 205100 71850
rect 204900 71620 205100 71650
rect 205400 71850 205600 71880
rect 205400 71650 205410 71850
rect 205480 71650 205520 71850
rect 205590 71650 205600 71850
rect 205400 71620 205600 71650
rect 205900 71850 206100 71880
rect 205900 71650 205910 71850
rect 205980 71650 206020 71850
rect 206090 71650 206100 71850
rect 205900 71620 206100 71650
rect 206400 71850 206600 71880
rect 206400 71650 206410 71850
rect 206480 71650 206520 71850
rect 206590 71650 206600 71850
rect 206400 71620 206600 71650
rect 206900 71850 207100 71880
rect 206900 71650 206910 71850
rect 206980 71650 207020 71850
rect 207090 71650 207100 71850
rect 206900 71620 207100 71650
rect 207400 71850 207600 71880
rect 207400 71650 207410 71850
rect 207480 71650 207520 71850
rect 207590 71650 207600 71850
rect 207400 71620 207600 71650
rect 207900 71850 208000 71880
rect 207900 71650 207910 71850
rect 207980 71650 208000 71850
rect 207900 71620 208000 71650
rect 196000 71600 196120 71620
rect 196380 71600 196620 71620
rect 196880 71600 197120 71620
rect 197380 71600 197620 71620
rect 197880 71600 198120 71620
rect 198380 71600 198620 71620
rect 198880 71600 199120 71620
rect 199380 71600 199620 71620
rect 199880 71600 200120 71620
rect 200380 71600 200620 71620
rect 200880 71600 201120 71620
rect 201380 71600 201620 71620
rect 201880 71600 202120 71620
rect 202380 71600 202620 71620
rect 202880 71600 203120 71620
rect 203380 71600 203620 71620
rect 203880 71600 204120 71620
rect 204380 71600 204620 71620
rect 204880 71600 205120 71620
rect 205380 71600 205620 71620
rect 205880 71600 206120 71620
rect 206380 71600 206620 71620
rect 206880 71600 207120 71620
rect 207380 71600 207620 71620
rect 207880 71600 208000 71620
rect 196000 71590 208000 71600
rect 196000 71520 196150 71590
rect 196350 71520 196650 71590
rect 196850 71520 197150 71590
rect 197350 71520 197650 71590
rect 197850 71520 198150 71590
rect 198350 71520 198650 71590
rect 198850 71520 199150 71590
rect 199350 71520 199650 71590
rect 199850 71520 200150 71590
rect 200350 71520 200650 71590
rect 200850 71520 201150 71590
rect 201350 71520 201650 71590
rect 201850 71520 202150 71590
rect 202350 71520 202650 71590
rect 202850 71520 203150 71590
rect 203350 71520 203650 71590
rect 203850 71520 204150 71590
rect 204350 71520 204650 71590
rect 204850 71520 205150 71590
rect 205350 71520 205650 71590
rect 205850 71520 206150 71590
rect 206350 71520 206650 71590
rect 206850 71520 207150 71590
rect 207350 71520 207650 71590
rect 207850 71520 208000 71590
rect 196000 71480 208000 71520
rect 196000 71410 196150 71480
rect 196350 71410 196650 71480
rect 196850 71410 197150 71480
rect 197350 71410 197650 71480
rect 197850 71410 198150 71480
rect 198350 71410 198650 71480
rect 198850 71410 199150 71480
rect 199350 71410 199650 71480
rect 199850 71410 200150 71480
rect 200350 71410 200650 71480
rect 200850 71410 201150 71480
rect 201350 71410 201650 71480
rect 201850 71410 202150 71480
rect 202350 71410 202650 71480
rect 202850 71410 203150 71480
rect 203350 71410 203650 71480
rect 203850 71410 204150 71480
rect 204350 71410 204650 71480
rect 204850 71410 205150 71480
rect 205350 71410 205650 71480
rect 205850 71410 206150 71480
rect 206350 71410 206650 71480
rect 206850 71410 207150 71480
rect 207350 71410 207650 71480
rect 207850 71410 208000 71480
rect 196000 71400 208000 71410
rect 196000 71380 196120 71400
rect 196380 71380 196620 71400
rect 196880 71380 197120 71400
rect 197380 71380 197620 71400
rect 197880 71380 198120 71400
rect 198380 71380 198620 71400
rect 198880 71380 199120 71400
rect 199380 71380 199620 71400
rect 199880 71380 200120 71400
rect 200380 71380 200620 71400
rect 200880 71380 201120 71400
rect 201380 71380 201620 71400
rect 201880 71380 202120 71400
rect 202380 71380 202620 71400
rect 202880 71380 203120 71400
rect 203380 71380 203620 71400
rect 203880 71380 204120 71400
rect 204380 71380 204620 71400
rect 204880 71380 205120 71400
rect 205380 71380 205620 71400
rect 205880 71380 206120 71400
rect 206380 71380 206620 71400
rect 206880 71380 207120 71400
rect 207380 71380 207620 71400
rect 207880 71380 208000 71400
rect 196000 71350 196100 71380
rect 196000 71150 196020 71350
rect 196090 71150 196100 71350
rect 196000 71120 196100 71150
rect 196400 71350 196600 71380
rect 196400 71150 196410 71350
rect 196480 71150 196520 71350
rect 196590 71150 196600 71350
rect 196400 71120 196600 71150
rect 196900 71350 197100 71380
rect 196900 71150 196910 71350
rect 196980 71150 197020 71350
rect 197090 71150 197100 71350
rect 196900 71120 197100 71150
rect 197400 71350 197600 71380
rect 197400 71150 197410 71350
rect 197480 71150 197520 71350
rect 197590 71150 197600 71350
rect 197400 71120 197600 71150
rect 197900 71350 198100 71380
rect 197900 71150 197910 71350
rect 197980 71150 198020 71350
rect 198090 71150 198100 71350
rect 197900 71120 198100 71150
rect 198400 71350 198600 71380
rect 198400 71150 198410 71350
rect 198480 71150 198520 71350
rect 198590 71150 198600 71350
rect 198400 71120 198600 71150
rect 198900 71350 199100 71380
rect 198900 71150 198910 71350
rect 198980 71150 199020 71350
rect 199090 71150 199100 71350
rect 198900 71120 199100 71150
rect 199400 71350 199600 71380
rect 199400 71150 199410 71350
rect 199480 71150 199520 71350
rect 199590 71150 199600 71350
rect 199400 71120 199600 71150
rect 199900 71350 200100 71380
rect 199900 71150 199910 71350
rect 199980 71150 200020 71350
rect 200090 71150 200100 71350
rect 199900 71120 200100 71150
rect 200400 71350 200600 71380
rect 200400 71150 200410 71350
rect 200480 71150 200520 71350
rect 200590 71150 200600 71350
rect 200400 71120 200600 71150
rect 200900 71350 201100 71380
rect 200900 71150 200910 71350
rect 200980 71150 201020 71350
rect 201090 71150 201100 71350
rect 200900 71120 201100 71150
rect 201400 71350 201600 71380
rect 201400 71150 201410 71350
rect 201480 71150 201520 71350
rect 201590 71150 201600 71350
rect 201400 71120 201600 71150
rect 201900 71350 202100 71380
rect 201900 71150 201910 71350
rect 201980 71150 202020 71350
rect 202090 71150 202100 71350
rect 201900 71120 202100 71150
rect 202400 71350 202600 71380
rect 202400 71150 202410 71350
rect 202480 71150 202520 71350
rect 202590 71150 202600 71350
rect 202400 71120 202600 71150
rect 202900 71350 203100 71380
rect 202900 71150 202910 71350
rect 202980 71150 203020 71350
rect 203090 71150 203100 71350
rect 202900 71120 203100 71150
rect 203400 71350 203600 71380
rect 203400 71150 203410 71350
rect 203480 71150 203520 71350
rect 203590 71150 203600 71350
rect 203400 71120 203600 71150
rect 203900 71350 204100 71380
rect 203900 71150 203910 71350
rect 203980 71150 204020 71350
rect 204090 71150 204100 71350
rect 203900 71120 204100 71150
rect 204400 71350 204600 71380
rect 204400 71150 204410 71350
rect 204480 71150 204520 71350
rect 204590 71150 204600 71350
rect 204400 71120 204600 71150
rect 204900 71350 205100 71380
rect 204900 71150 204910 71350
rect 204980 71150 205020 71350
rect 205090 71150 205100 71350
rect 204900 71120 205100 71150
rect 205400 71350 205600 71380
rect 205400 71150 205410 71350
rect 205480 71150 205520 71350
rect 205590 71150 205600 71350
rect 205400 71120 205600 71150
rect 205900 71350 206100 71380
rect 205900 71150 205910 71350
rect 205980 71150 206020 71350
rect 206090 71150 206100 71350
rect 205900 71120 206100 71150
rect 206400 71350 206600 71380
rect 206400 71150 206410 71350
rect 206480 71150 206520 71350
rect 206590 71150 206600 71350
rect 206400 71120 206600 71150
rect 206900 71350 207100 71380
rect 206900 71150 206910 71350
rect 206980 71150 207020 71350
rect 207090 71150 207100 71350
rect 206900 71120 207100 71150
rect 207400 71350 207600 71380
rect 207400 71150 207410 71350
rect 207480 71150 207520 71350
rect 207590 71150 207600 71350
rect 207400 71120 207600 71150
rect 207900 71350 208000 71380
rect 207900 71150 207910 71350
rect 207980 71150 208000 71350
rect 207900 71120 208000 71150
rect 196000 71100 196120 71120
rect 196380 71100 196620 71120
rect 196880 71100 197120 71120
rect 197380 71100 197620 71120
rect 197880 71100 198120 71120
rect 198380 71100 198620 71120
rect 198880 71100 199120 71120
rect 199380 71100 199620 71120
rect 199880 71100 200120 71120
rect 200380 71100 200620 71120
rect 200880 71100 201120 71120
rect 201380 71100 201620 71120
rect 201880 71100 202120 71120
rect 202380 71100 202620 71120
rect 202880 71100 203120 71120
rect 203380 71100 203620 71120
rect 203880 71100 204120 71120
rect 204380 71100 204620 71120
rect 204880 71100 205120 71120
rect 205380 71100 205620 71120
rect 205880 71100 206120 71120
rect 206380 71100 206620 71120
rect 206880 71100 207120 71120
rect 207380 71100 207620 71120
rect 207880 71100 208000 71120
rect 196000 71090 208000 71100
rect 196000 71020 196150 71090
rect 196350 71020 196650 71090
rect 196850 71020 197150 71090
rect 197350 71020 197650 71090
rect 197850 71020 198150 71090
rect 198350 71020 198650 71090
rect 198850 71020 199150 71090
rect 199350 71020 199650 71090
rect 199850 71020 200150 71090
rect 200350 71020 200650 71090
rect 200850 71020 201150 71090
rect 201350 71020 201650 71090
rect 201850 71020 202150 71090
rect 202350 71020 202650 71090
rect 202850 71020 203150 71090
rect 203350 71020 203650 71090
rect 203850 71020 204150 71090
rect 204350 71020 204650 71090
rect 204850 71020 205150 71090
rect 205350 71020 205650 71090
rect 205850 71020 206150 71090
rect 206350 71020 206650 71090
rect 206850 71020 207150 71090
rect 207350 71020 207650 71090
rect 207850 71020 208000 71090
rect 196000 70980 208000 71020
rect 196000 70910 196150 70980
rect 196350 70910 196650 70980
rect 196850 70910 197150 70980
rect 197350 70910 197650 70980
rect 197850 70910 198150 70980
rect 198350 70910 198650 70980
rect 198850 70910 199150 70980
rect 199350 70910 199650 70980
rect 199850 70910 200150 70980
rect 200350 70910 200650 70980
rect 200850 70910 201150 70980
rect 201350 70910 201650 70980
rect 201850 70910 202150 70980
rect 202350 70910 202650 70980
rect 202850 70910 203150 70980
rect 203350 70910 203650 70980
rect 203850 70910 204150 70980
rect 204350 70910 204650 70980
rect 204850 70910 205150 70980
rect 205350 70910 205650 70980
rect 205850 70910 206150 70980
rect 206350 70910 206650 70980
rect 206850 70910 207150 70980
rect 207350 70910 207650 70980
rect 207850 70910 208000 70980
rect 196000 70900 208000 70910
rect 196000 70880 196120 70900
rect 196380 70880 196620 70900
rect 196880 70880 197120 70900
rect 197380 70880 197620 70900
rect 197880 70880 198120 70900
rect 198380 70880 198620 70900
rect 198880 70880 199120 70900
rect 199380 70880 199620 70900
rect 199880 70880 200120 70900
rect 200380 70880 200620 70900
rect 200880 70880 201120 70900
rect 201380 70880 201620 70900
rect 201880 70880 202120 70900
rect 202380 70880 202620 70900
rect 202880 70880 203120 70900
rect 203380 70880 203620 70900
rect 203880 70880 204120 70900
rect 204380 70880 204620 70900
rect 204880 70880 205120 70900
rect 205380 70880 205620 70900
rect 205880 70880 206120 70900
rect 206380 70880 206620 70900
rect 206880 70880 207120 70900
rect 207380 70880 207620 70900
rect 207880 70880 208000 70900
rect 196000 70850 196100 70880
rect 196000 70650 196020 70850
rect 196090 70650 196100 70850
rect 196000 70620 196100 70650
rect 196400 70850 196600 70880
rect 196400 70650 196410 70850
rect 196480 70650 196520 70850
rect 196590 70650 196600 70850
rect 196400 70620 196600 70650
rect 196900 70850 197100 70880
rect 196900 70650 196910 70850
rect 196980 70650 197020 70850
rect 197090 70650 197100 70850
rect 196900 70620 197100 70650
rect 197400 70850 197600 70880
rect 197400 70650 197410 70850
rect 197480 70650 197520 70850
rect 197590 70650 197600 70850
rect 197400 70620 197600 70650
rect 197900 70850 198100 70880
rect 197900 70650 197910 70850
rect 197980 70650 198020 70850
rect 198090 70650 198100 70850
rect 197900 70620 198100 70650
rect 198400 70850 198600 70880
rect 198400 70650 198410 70850
rect 198480 70650 198520 70850
rect 198590 70650 198600 70850
rect 198400 70620 198600 70650
rect 198900 70850 199100 70880
rect 198900 70650 198910 70850
rect 198980 70650 199020 70850
rect 199090 70650 199100 70850
rect 198900 70620 199100 70650
rect 199400 70850 199600 70880
rect 199400 70650 199410 70850
rect 199480 70650 199520 70850
rect 199590 70650 199600 70850
rect 199400 70620 199600 70650
rect 199900 70850 200100 70880
rect 199900 70650 199910 70850
rect 199980 70650 200020 70850
rect 200090 70650 200100 70850
rect 199900 70620 200100 70650
rect 200400 70850 200600 70880
rect 200400 70650 200410 70850
rect 200480 70650 200520 70850
rect 200590 70650 200600 70850
rect 200400 70620 200600 70650
rect 200900 70850 201100 70880
rect 200900 70650 200910 70850
rect 200980 70650 201020 70850
rect 201090 70650 201100 70850
rect 200900 70620 201100 70650
rect 201400 70850 201600 70880
rect 201400 70650 201410 70850
rect 201480 70650 201520 70850
rect 201590 70650 201600 70850
rect 201400 70620 201600 70650
rect 201900 70850 202100 70880
rect 201900 70650 201910 70850
rect 201980 70650 202020 70850
rect 202090 70650 202100 70850
rect 201900 70620 202100 70650
rect 202400 70850 202600 70880
rect 202400 70650 202410 70850
rect 202480 70650 202520 70850
rect 202590 70650 202600 70850
rect 202400 70620 202600 70650
rect 202900 70850 203100 70880
rect 202900 70650 202910 70850
rect 202980 70650 203020 70850
rect 203090 70650 203100 70850
rect 202900 70620 203100 70650
rect 203400 70850 203600 70880
rect 203400 70650 203410 70850
rect 203480 70650 203520 70850
rect 203590 70650 203600 70850
rect 203400 70620 203600 70650
rect 203900 70850 204100 70880
rect 203900 70650 203910 70850
rect 203980 70650 204020 70850
rect 204090 70650 204100 70850
rect 203900 70620 204100 70650
rect 204400 70850 204600 70880
rect 204400 70650 204410 70850
rect 204480 70650 204520 70850
rect 204590 70650 204600 70850
rect 204400 70620 204600 70650
rect 204900 70850 205100 70880
rect 204900 70650 204910 70850
rect 204980 70650 205020 70850
rect 205090 70650 205100 70850
rect 204900 70620 205100 70650
rect 205400 70850 205600 70880
rect 205400 70650 205410 70850
rect 205480 70650 205520 70850
rect 205590 70650 205600 70850
rect 205400 70620 205600 70650
rect 205900 70850 206100 70880
rect 205900 70650 205910 70850
rect 205980 70650 206020 70850
rect 206090 70650 206100 70850
rect 205900 70620 206100 70650
rect 206400 70850 206600 70880
rect 206400 70650 206410 70850
rect 206480 70650 206520 70850
rect 206590 70650 206600 70850
rect 206400 70620 206600 70650
rect 206900 70850 207100 70880
rect 206900 70650 206910 70850
rect 206980 70650 207020 70850
rect 207090 70650 207100 70850
rect 206900 70620 207100 70650
rect 207400 70850 207600 70880
rect 207400 70650 207410 70850
rect 207480 70650 207520 70850
rect 207590 70650 207600 70850
rect 207400 70620 207600 70650
rect 207900 70850 208000 70880
rect 207900 70650 207910 70850
rect 207980 70650 208000 70850
rect 207900 70620 208000 70650
rect 196000 70600 196120 70620
rect 196380 70600 196620 70620
rect 196880 70600 197120 70620
rect 197380 70600 197620 70620
rect 197880 70600 198120 70620
rect 198380 70600 198620 70620
rect 198880 70600 199120 70620
rect 199380 70600 199620 70620
rect 199880 70600 200120 70620
rect 200380 70600 200620 70620
rect 200880 70600 201120 70620
rect 201380 70600 201620 70620
rect 201880 70600 202120 70620
rect 202380 70600 202620 70620
rect 202880 70600 203120 70620
rect 203380 70600 203620 70620
rect 203880 70600 204120 70620
rect 204380 70600 204620 70620
rect 204880 70600 205120 70620
rect 205380 70600 205620 70620
rect 205880 70600 206120 70620
rect 206380 70600 206620 70620
rect 206880 70600 207120 70620
rect 207380 70600 207620 70620
rect 207880 70600 208000 70620
rect 196000 70590 208000 70600
rect 196000 70520 196150 70590
rect 196350 70520 196650 70590
rect 196850 70520 197150 70590
rect 197350 70520 197650 70590
rect 197850 70520 198150 70590
rect 198350 70520 198650 70590
rect 198850 70520 199150 70590
rect 199350 70520 199650 70590
rect 199850 70520 200150 70590
rect 200350 70520 200650 70590
rect 200850 70520 201150 70590
rect 201350 70520 201650 70590
rect 201850 70520 202150 70590
rect 202350 70520 202650 70590
rect 202850 70520 203150 70590
rect 203350 70520 203650 70590
rect 203850 70520 204150 70590
rect 204350 70520 204650 70590
rect 204850 70520 205150 70590
rect 205350 70520 205650 70590
rect 205850 70520 206150 70590
rect 206350 70520 206650 70590
rect 206850 70520 207150 70590
rect 207350 70520 207650 70590
rect 207850 70520 208000 70590
rect 196000 70480 208000 70520
rect 196000 70410 196150 70480
rect 196350 70410 196650 70480
rect 196850 70410 197150 70480
rect 197350 70410 197650 70480
rect 197850 70410 198150 70480
rect 198350 70410 198650 70480
rect 198850 70410 199150 70480
rect 199350 70410 199650 70480
rect 199850 70410 200150 70480
rect 200350 70410 200650 70480
rect 200850 70410 201150 70480
rect 201350 70410 201650 70480
rect 201850 70410 202150 70480
rect 202350 70410 202650 70480
rect 202850 70410 203150 70480
rect 203350 70410 203650 70480
rect 203850 70410 204150 70480
rect 204350 70410 204650 70480
rect 204850 70410 205150 70480
rect 205350 70410 205650 70480
rect 205850 70410 206150 70480
rect 206350 70410 206650 70480
rect 206850 70410 207150 70480
rect 207350 70410 207650 70480
rect 207850 70410 208000 70480
rect 196000 70400 208000 70410
rect 196000 70380 196120 70400
rect 196380 70380 196620 70400
rect 196880 70380 197120 70400
rect 197380 70380 197620 70400
rect 197880 70380 198120 70400
rect 198380 70380 198620 70400
rect 198880 70380 199120 70400
rect 199380 70380 199620 70400
rect 199880 70380 200120 70400
rect 200380 70380 200620 70400
rect 200880 70380 201120 70400
rect 201380 70380 201620 70400
rect 201880 70380 202120 70400
rect 202380 70380 202620 70400
rect 202880 70380 203120 70400
rect 203380 70380 203620 70400
rect 203880 70380 204120 70400
rect 204380 70380 204620 70400
rect 204880 70380 205120 70400
rect 205380 70380 205620 70400
rect 205880 70380 206120 70400
rect 206380 70380 206620 70400
rect 206880 70380 207120 70400
rect 207380 70380 207620 70400
rect 207880 70380 208000 70400
rect 196000 70350 196100 70380
rect 196000 70150 196020 70350
rect 196090 70150 196100 70350
rect 196000 70120 196100 70150
rect 196400 70350 196600 70380
rect 196400 70150 196410 70350
rect 196480 70150 196520 70350
rect 196590 70150 196600 70350
rect 196400 70120 196600 70150
rect 196900 70350 197100 70380
rect 196900 70150 196910 70350
rect 196980 70150 197020 70350
rect 197090 70150 197100 70350
rect 196900 70120 197100 70150
rect 197400 70350 197600 70380
rect 197400 70150 197410 70350
rect 197480 70150 197520 70350
rect 197590 70150 197600 70350
rect 197400 70120 197600 70150
rect 197900 70350 198100 70380
rect 197900 70150 197910 70350
rect 197980 70150 198020 70350
rect 198090 70150 198100 70350
rect 197900 70120 198100 70150
rect 198400 70350 198600 70380
rect 198400 70150 198410 70350
rect 198480 70150 198520 70350
rect 198590 70150 198600 70350
rect 198400 70120 198600 70150
rect 198900 70350 199100 70380
rect 198900 70150 198910 70350
rect 198980 70150 199020 70350
rect 199090 70150 199100 70350
rect 198900 70120 199100 70150
rect 199400 70350 199600 70380
rect 199400 70150 199410 70350
rect 199480 70150 199520 70350
rect 199590 70150 199600 70350
rect 199400 70120 199600 70150
rect 199900 70350 200100 70380
rect 199900 70150 199910 70350
rect 199980 70150 200020 70350
rect 200090 70150 200100 70350
rect 199900 70120 200100 70150
rect 200400 70350 200600 70380
rect 200400 70150 200410 70350
rect 200480 70150 200520 70350
rect 200590 70150 200600 70350
rect 200400 70120 200600 70150
rect 200900 70350 201100 70380
rect 200900 70150 200910 70350
rect 200980 70150 201020 70350
rect 201090 70150 201100 70350
rect 200900 70120 201100 70150
rect 201400 70350 201600 70380
rect 201400 70150 201410 70350
rect 201480 70150 201520 70350
rect 201590 70150 201600 70350
rect 201400 70120 201600 70150
rect 201900 70350 202100 70380
rect 201900 70150 201910 70350
rect 201980 70150 202020 70350
rect 202090 70150 202100 70350
rect 201900 70120 202100 70150
rect 202400 70350 202600 70380
rect 202400 70150 202410 70350
rect 202480 70150 202520 70350
rect 202590 70150 202600 70350
rect 202400 70120 202600 70150
rect 202900 70350 203100 70380
rect 202900 70150 202910 70350
rect 202980 70150 203020 70350
rect 203090 70150 203100 70350
rect 202900 70120 203100 70150
rect 203400 70350 203600 70380
rect 203400 70150 203410 70350
rect 203480 70150 203520 70350
rect 203590 70150 203600 70350
rect 203400 70120 203600 70150
rect 203900 70350 204100 70380
rect 203900 70150 203910 70350
rect 203980 70150 204020 70350
rect 204090 70150 204100 70350
rect 203900 70120 204100 70150
rect 204400 70350 204600 70380
rect 204400 70150 204410 70350
rect 204480 70150 204520 70350
rect 204590 70150 204600 70350
rect 204400 70120 204600 70150
rect 204900 70350 205100 70380
rect 204900 70150 204910 70350
rect 204980 70150 205020 70350
rect 205090 70150 205100 70350
rect 204900 70120 205100 70150
rect 205400 70350 205600 70380
rect 205400 70150 205410 70350
rect 205480 70150 205520 70350
rect 205590 70150 205600 70350
rect 205400 70120 205600 70150
rect 205900 70350 206100 70380
rect 205900 70150 205910 70350
rect 205980 70150 206020 70350
rect 206090 70150 206100 70350
rect 205900 70120 206100 70150
rect 206400 70350 206600 70380
rect 206400 70150 206410 70350
rect 206480 70150 206520 70350
rect 206590 70150 206600 70350
rect 206400 70120 206600 70150
rect 206900 70350 207100 70380
rect 206900 70150 206910 70350
rect 206980 70150 207020 70350
rect 207090 70150 207100 70350
rect 206900 70120 207100 70150
rect 207400 70350 207600 70380
rect 207400 70150 207410 70350
rect 207480 70150 207520 70350
rect 207590 70150 207600 70350
rect 207400 70120 207600 70150
rect 207900 70350 208000 70380
rect 207900 70150 207910 70350
rect 207980 70150 208000 70350
rect 207900 70120 208000 70150
rect 196000 70100 196120 70120
rect 196380 70100 196620 70120
rect 196880 70100 197120 70120
rect 197380 70100 197620 70120
rect 197880 70100 198120 70120
rect 198380 70100 198620 70120
rect 198880 70100 199120 70120
rect 199380 70100 199620 70120
rect 199880 70100 200120 70120
rect 200380 70100 200620 70120
rect 200880 70100 201120 70120
rect 201380 70100 201620 70120
rect 201880 70100 202120 70120
rect 202380 70100 202620 70120
rect 202880 70100 203120 70120
rect 203380 70100 203620 70120
rect 203880 70100 204120 70120
rect 204380 70100 204620 70120
rect 204880 70100 205120 70120
rect 205380 70100 205620 70120
rect 205880 70100 206120 70120
rect 206380 70100 206620 70120
rect 206880 70100 207120 70120
rect 207380 70100 207620 70120
rect 207880 70100 208000 70120
rect 196000 70090 208000 70100
rect 196000 70020 196150 70090
rect 196350 70020 196650 70090
rect 196850 70020 197150 70090
rect 197350 70020 197650 70090
rect 197850 70020 198150 70090
rect 198350 70020 198650 70090
rect 198850 70020 199150 70090
rect 199350 70020 199650 70090
rect 199850 70020 200150 70090
rect 200350 70020 200650 70090
rect 200850 70020 201150 70090
rect 201350 70020 201650 70090
rect 201850 70020 202150 70090
rect 202350 70020 202650 70090
rect 202850 70020 203150 70090
rect 203350 70020 203650 70090
rect 203850 70020 204150 70090
rect 204350 70020 204650 70090
rect 204850 70020 205150 70090
rect 205350 70020 205650 70090
rect 205850 70020 206150 70090
rect 206350 70020 206650 70090
rect 206850 70020 207150 70090
rect 207350 70020 207650 70090
rect 207850 70020 208000 70090
rect 196000 69980 208000 70020
rect 196000 69910 196150 69980
rect 196350 69910 196650 69980
rect 196850 69910 197150 69980
rect 197350 69910 197650 69980
rect 197850 69910 198150 69980
rect 198350 69910 198650 69980
rect 198850 69910 199150 69980
rect 199350 69910 199650 69980
rect 199850 69910 200150 69980
rect 200350 69910 200650 69980
rect 200850 69910 201150 69980
rect 201350 69910 201650 69980
rect 201850 69910 202150 69980
rect 202350 69910 202650 69980
rect 202850 69910 203150 69980
rect 203350 69910 203650 69980
rect 203850 69910 204150 69980
rect 204350 69910 204650 69980
rect 204850 69910 205150 69980
rect 205350 69910 205650 69980
rect 205850 69910 206150 69980
rect 206350 69910 206650 69980
rect 206850 69910 207150 69980
rect 207350 69910 207650 69980
rect 207850 69910 208000 69980
rect 196000 69900 208000 69910
rect 196000 69880 196120 69900
rect 196380 69880 196620 69900
rect 196880 69880 197120 69900
rect 197380 69880 197620 69900
rect 197880 69880 198120 69900
rect 198380 69880 198620 69900
rect 198880 69880 199120 69900
rect 199380 69880 199620 69900
rect 199880 69880 200120 69900
rect 200380 69880 200620 69900
rect 200880 69880 201120 69900
rect 201380 69880 201620 69900
rect 201880 69880 202120 69900
rect 202380 69880 202620 69900
rect 202880 69880 203120 69900
rect 203380 69880 203620 69900
rect 203880 69880 204120 69900
rect 204380 69880 204620 69900
rect 204880 69880 205120 69900
rect 205380 69880 205620 69900
rect 205880 69880 206120 69900
rect 206380 69880 206620 69900
rect 206880 69880 207120 69900
rect 207380 69880 207620 69900
rect 207880 69880 208000 69900
rect 196000 69850 196100 69880
rect 196000 69650 196020 69850
rect 196090 69650 196100 69850
rect 196000 69620 196100 69650
rect 196400 69850 196600 69880
rect 196400 69650 196410 69850
rect 196480 69650 196520 69850
rect 196590 69650 196600 69850
rect 196400 69620 196600 69650
rect 196900 69850 197100 69880
rect 196900 69650 196910 69850
rect 196980 69650 197020 69850
rect 197090 69650 197100 69850
rect 196900 69620 197100 69650
rect 197400 69850 197600 69880
rect 197400 69650 197410 69850
rect 197480 69650 197520 69850
rect 197590 69650 197600 69850
rect 197400 69620 197600 69650
rect 197900 69850 198100 69880
rect 197900 69650 197910 69850
rect 197980 69650 198020 69850
rect 198090 69650 198100 69850
rect 197900 69620 198100 69650
rect 198400 69850 198600 69880
rect 198400 69650 198410 69850
rect 198480 69650 198520 69850
rect 198590 69650 198600 69850
rect 198400 69620 198600 69650
rect 198900 69850 199100 69880
rect 198900 69650 198910 69850
rect 198980 69650 199020 69850
rect 199090 69650 199100 69850
rect 198900 69620 199100 69650
rect 199400 69850 199600 69880
rect 199400 69650 199410 69850
rect 199480 69650 199520 69850
rect 199590 69650 199600 69850
rect 199400 69620 199600 69650
rect 199900 69850 200100 69880
rect 199900 69650 199910 69850
rect 199980 69650 200020 69850
rect 200090 69650 200100 69850
rect 199900 69620 200100 69650
rect 200400 69850 200600 69880
rect 200400 69650 200410 69850
rect 200480 69650 200520 69850
rect 200590 69650 200600 69850
rect 200400 69620 200600 69650
rect 200900 69850 201100 69880
rect 200900 69650 200910 69850
rect 200980 69650 201020 69850
rect 201090 69650 201100 69850
rect 200900 69620 201100 69650
rect 201400 69850 201600 69880
rect 201400 69650 201410 69850
rect 201480 69650 201520 69850
rect 201590 69650 201600 69850
rect 201400 69620 201600 69650
rect 201900 69850 202100 69880
rect 201900 69650 201910 69850
rect 201980 69650 202020 69850
rect 202090 69650 202100 69850
rect 201900 69620 202100 69650
rect 202400 69850 202600 69880
rect 202400 69650 202410 69850
rect 202480 69650 202520 69850
rect 202590 69650 202600 69850
rect 202400 69620 202600 69650
rect 202900 69850 203100 69880
rect 202900 69650 202910 69850
rect 202980 69650 203020 69850
rect 203090 69650 203100 69850
rect 202900 69620 203100 69650
rect 203400 69850 203600 69880
rect 203400 69650 203410 69850
rect 203480 69650 203520 69850
rect 203590 69650 203600 69850
rect 203400 69620 203600 69650
rect 203900 69850 204100 69880
rect 203900 69650 203910 69850
rect 203980 69650 204020 69850
rect 204090 69650 204100 69850
rect 203900 69620 204100 69650
rect 204400 69850 204600 69880
rect 204400 69650 204410 69850
rect 204480 69650 204520 69850
rect 204590 69650 204600 69850
rect 204400 69620 204600 69650
rect 204900 69850 205100 69880
rect 204900 69650 204910 69850
rect 204980 69650 205020 69850
rect 205090 69650 205100 69850
rect 204900 69620 205100 69650
rect 205400 69850 205600 69880
rect 205400 69650 205410 69850
rect 205480 69650 205520 69850
rect 205590 69650 205600 69850
rect 205400 69620 205600 69650
rect 205900 69850 206100 69880
rect 205900 69650 205910 69850
rect 205980 69650 206020 69850
rect 206090 69650 206100 69850
rect 205900 69620 206100 69650
rect 206400 69850 206600 69880
rect 206400 69650 206410 69850
rect 206480 69650 206520 69850
rect 206590 69650 206600 69850
rect 206400 69620 206600 69650
rect 206900 69850 207100 69880
rect 206900 69650 206910 69850
rect 206980 69650 207020 69850
rect 207090 69650 207100 69850
rect 206900 69620 207100 69650
rect 207400 69850 207600 69880
rect 207400 69650 207410 69850
rect 207480 69650 207520 69850
rect 207590 69650 207600 69850
rect 207400 69620 207600 69650
rect 207900 69850 208000 69880
rect 207900 69650 207910 69850
rect 207980 69650 208000 69850
rect 207900 69620 208000 69650
rect 196000 69600 196120 69620
rect 196380 69600 196620 69620
rect 196880 69600 197120 69620
rect 197380 69600 197620 69620
rect 197880 69600 198120 69620
rect 198380 69600 198620 69620
rect 198880 69600 199120 69620
rect 199380 69600 199620 69620
rect 199880 69600 200120 69620
rect 200380 69600 200620 69620
rect 200880 69600 201120 69620
rect 201380 69600 201620 69620
rect 201880 69600 202120 69620
rect 202380 69600 202620 69620
rect 202880 69600 203120 69620
rect 203380 69600 203620 69620
rect 203880 69600 204120 69620
rect 204380 69600 204620 69620
rect 204880 69600 205120 69620
rect 205380 69600 205620 69620
rect 205880 69600 206120 69620
rect 206380 69600 206620 69620
rect 206880 69600 207120 69620
rect 207380 69600 207620 69620
rect 207880 69600 208000 69620
rect 196000 69590 208000 69600
rect 196000 69520 196150 69590
rect 196350 69520 196650 69590
rect 196850 69520 197150 69590
rect 197350 69520 197650 69590
rect 197850 69520 198150 69590
rect 198350 69520 198650 69590
rect 198850 69520 199150 69590
rect 199350 69520 199650 69590
rect 199850 69520 200150 69590
rect 200350 69520 200650 69590
rect 200850 69520 201150 69590
rect 201350 69520 201650 69590
rect 201850 69520 202150 69590
rect 202350 69520 202650 69590
rect 202850 69520 203150 69590
rect 203350 69520 203650 69590
rect 203850 69520 204150 69590
rect 204350 69520 204650 69590
rect 204850 69520 205150 69590
rect 205350 69520 205650 69590
rect 205850 69520 206150 69590
rect 206350 69520 206650 69590
rect 206850 69520 207150 69590
rect 207350 69520 207650 69590
rect 207850 69520 208000 69590
rect 196000 69480 208000 69520
rect 196000 69410 196150 69480
rect 196350 69410 196650 69480
rect 196850 69410 197150 69480
rect 197350 69410 197650 69480
rect 197850 69410 198150 69480
rect 198350 69410 198650 69480
rect 198850 69410 199150 69480
rect 199350 69410 199650 69480
rect 199850 69410 200150 69480
rect 200350 69410 200650 69480
rect 200850 69410 201150 69480
rect 201350 69410 201650 69480
rect 201850 69410 202150 69480
rect 202350 69410 202650 69480
rect 202850 69410 203150 69480
rect 203350 69410 203650 69480
rect 203850 69410 204150 69480
rect 204350 69410 204650 69480
rect 204850 69410 205150 69480
rect 205350 69410 205650 69480
rect 205850 69410 206150 69480
rect 206350 69410 206650 69480
rect 206850 69410 207150 69480
rect 207350 69410 207650 69480
rect 207850 69410 208000 69480
rect 196000 69400 208000 69410
rect 196000 69380 196120 69400
rect 196380 69380 196620 69400
rect 196880 69380 197120 69400
rect 197380 69380 197620 69400
rect 197880 69380 198120 69400
rect 198380 69380 198620 69400
rect 198880 69380 199120 69400
rect 199380 69380 199620 69400
rect 199880 69380 200120 69400
rect 200380 69380 200620 69400
rect 200880 69380 201120 69400
rect 201380 69380 201620 69400
rect 201880 69380 202120 69400
rect 202380 69380 202620 69400
rect 202880 69380 203120 69400
rect 203380 69380 203620 69400
rect 203880 69380 204120 69400
rect 204380 69380 204620 69400
rect 204880 69380 205120 69400
rect 205380 69380 205620 69400
rect 205880 69380 206120 69400
rect 206380 69380 206620 69400
rect 206880 69380 207120 69400
rect 207380 69380 207620 69400
rect 207880 69380 208000 69400
rect 196000 69350 196100 69380
rect 196000 69150 196020 69350
rect 196090 69150 196100 69350
rect 196000 69120 196100 69150
rect 196400 69350 196600 69380
rect 196400 69150 196410 69350
rect 196480 69150 196520 69350
rect 196590 69150 196600 69350
rect 196400 69120 196600 69150
rect 196900 69350 197100 69380
rect 196900 69150 196910 69350
rect 196980 69150 197020 69350
rect 197090 69150 197100 69350
rect 196900 69120 197100 69150
rect 197400 69350 197600 69380
rect 197400 69150 197410 69350
rect 197480 69150 197520 69350
rect 197590 69150 197600 69350
rect 197400 69120 197600 69150
rect 197900 69350 198100 69380
rect 197900 69150 197910 69350
rect 197980 69150 198020 69350
rect 198090 69150 198100 69350
rect 197900 69120 198100 69150
rect 198400 69350 198600 69380
rect 198400 69150 198410 69350
rect 198480 69150 198520 69350
rect 198590 69150 198600 69350
rect 198400 69120 198600 69150
rect 198900 69350 199100 69380
rect 198900 69150 198910 69350
rect 198980 69150 199020 69350
rect 199090 69150 199100 69350
rect 198900 69120 199100 69150
rect 199400 69350 199600 69380
rect 199400 69150 199410 69350
rect 199480 69150 199520 69350
rect 199590 69150 199600 69350
rect 199400 69120 199600 69150
rect 199900 69350 200100 69380
rect 199900 69150 199910 69350
rect 199980 69150 200020 69350
rect 200090 69150 200100 69350
rect 199900 69120 200100 69150
rect 200400 69350 200600 69380
rect 200400 69150 200410 69350
rect 200480 69150 200520 69350
rect 200590 69150 200600 69350
rect 200400 69120 200600 69150
rect 200900 69350 201100 69380
rect 200900 69150 200910 69350
rect 200980 69150 201020 69350
rect 201090 69150 201100 69350
rect 200900 69120 201100 69150
rect 201400 69350 201600 69380
rect 201400 69150 201410 69350
rect 201480 69150 201520 69350
rect 201590 69150 201600 69350
rect 201400 69120 201600 69150
rect 201900 69350 202100 69380
rect 201900 69150 201910 69350
rect 201980 69150 202020 69350
rect 202090 69150 202100 69350
rect 201900 69120 202100 69150
rect 202400 69350 202600 69380
rect 202400 69150 202410 69350
rect 202480 69150 202520 69350
rect 202590 69150 202600 69350
rect 202400 69120 202600 69150
rect 202900 69350 203100 69380
rect 202900 69150 202910 69350
rect 202980 69150 203020 69350
rect 203090 69150 203100 69350
rect 202900 69120 203100 69150
rect 203400 69350 203600 69380
rect 203400 69150 203410 69350
rect 203480 69150 203520 69350
rect 203590 69150 203600 69350
rect 203400 69120 203600 69150
rect 203900 69350 204100 69380
rect 203900 69150 203910 69350
rect 203980 69150 204020 69350
rect 204090 69150 204100 69350
rect 203900 69120 204100 69150
rect 204400 69350 204600 69380
rect 204400 69150 204410 69350
rect 204480 69150 204520 69350
rect 204590 69150 204600 69350
rect 204400 69120 204600 69150
rect 204900 69350 205100 69380
rect 204900 69150 204910 69350
rect 204980 69150 205020 69350
rect 205090 69150 205100 69350
rect 204900 69120 205100 69150
rect 205400 69350 205600 69380
rect 205400 69150 205410 69350
rect 205480 69150 205520 69350
rect 205590 69150 205600 69350
rect 205400 69120 205600 69150
rect 205900 69350 206100 69380
rect 205900 69150 205910 69350
rect 205980 69150 206020 69350
rect 206090 69150 206100 69350
rect 205900 69120 206100 69150
rect 206400 69350 206600 69380
rect 206400 69150 206410 69350
rect 206480 69150 206520 69350
rect 206590 69150 206600 69350
rect 206400 69120 206600 69150
rect 206900 69350 207100 69380
rect 206900 69150 206910 69350
rect 206980 69150 207020 69350
rect 207090 69150 207100 69350
rect 206900 69120 207100 69150
rect 207400 69350 207600 69380
rect 207400 69150 207410 69350
rect 207480 69150 207520 69350
rect 207590 69150 207600 69350
rect 207400 69120 207600 69150
rect 207900 69350 208000 69380
rect 207900 69150 207910 69350
rect 207980 69150 208000 69350
rect 207900 69120 208000 69150
rect 196000 69100 196120 69120
rect 196380 69100 196620 69120
rect 196880 69100 197120 69120
rect 197380 69100 197620 69120
rect 197880 69100 198120 69120
rect 198380 69100 198620 69120
rect 198880 69100 199120 69120
rect 199380 69100 199620 69120
rect 199880 69100 200120 69120
rect 200380 69100 200620 69120
rect 200880 69100 201120 69120
rect 201380 69100 201620 69120
rect 201880 69100 202120 69120
rect 202380 69100 202620 69120
rect 202880 69100 203120 69120
rect 203380 69100 203620 69120
rect 203880 69100 204120 69120
rect 204380 69100 204620 69120
rect 204880 69100 205120 69120
rect 205380 69100 205620 69120
rect 205880 69100 206120 69120
rect 206380 69100 206620 69120
rect 206880 69100 207120 69120
rect 207380 69100 207620 69120
rect 207880 69100 208000 69120
rect 196000 69090 208000 69100
rect 196000 69020 196150 69090
rect 196350 69020 196650 69090
rect 196850 69020 197150 69090
rect 197350 69020 197650 69090
rect 197850 69020 198150 69090
rect 198350 69020 198650 69090
rect 198850 69020 199150 69090
rect 199350 69020 199650 69090
rect 199850 69020 200150 69090
rect 200350 69020 200650 69090
rect 200850 69020 201150 69090
rect 201350 69020 201650 69090
rect 201850 69020 202150 69090
rect 202350 69020 202650 69090
rect 202850 69020 203150 69090
rect 203350 69020 203650 69090
rect 203850 69020 204150 69090
rect 204350 69020 204650 69090
rect 204850 69020 205150 69090
rect 205350 69020 205650 69090
rect 205850 69020 206150 69090
rect 206350 69020 206650 69090
rect 206850 69020 207150 69090
rect 207350 69020 207650 69090
rect 207850 69020 208000 69090
rect 196000 68980 208000 69020
rect 196000 68910 196150 68980
rect 196350 68910 196650 68980
rect 196850 68910 197150 68980
rect 197350 68910 197650 68980
rect 197850 68910 198150 68980
rect 198350 68910 198650 68980
rect 198850 68910 199150 68980
rect 199350 68910 199650 68980
rect 199850 68910 200150 68980
rect 200350 68910 200650 68980
rect 200850 68910 201150 68980
rect 201350 68910 201650 68980
rect 201850 68910 202150 68980
rect 202350 68910 202650 68980
rect 202850 68910 203150 68980
rect 203350 68910 203650 68980
rect 203850 68910 204150 68980
rect 204350 68910 204650 68980
rect 204850 68910 205150 68980
rect 205350 68910 205650 68980
rect 205850 68910 206150 68980
rect 206350 68910 206650 68980
rect 206850 68910 207150 68980
rect 207350 68910 207650 68980
rect 207850 68910 208000 68980
rect 196000 68900 208000 68910
rect 196000 68880 196120 68900
rect 196380 68880 196620 68900
rect 196880 68880 197120 68900
rect 197380 68880 197620 68900
rect 197880 68880 198120 68900
rect 198380 68880 198620 68900
rect 198880 68880 199120 68900
rect 199380 68880 199620 68900
rect 199880 68880 200120 68900
rect 200380 68880 200620 68900
rect 200880 68880 201120 68900
rect 201380 68880 201620 68900
rect 201880 68880 202120 68900
rect 202380 68880 202620 68900
rect 202880 68880 203120 68900
rect 203380 68880 203620 68900
rect 203880 68880 204120 68900
rect 204380 68880 204620 68900
rect 204880 68880 205120 68900
rect 205380 68880 205620 68900
rect 205880 68880 206120 68900
rect 206380 68880 206620 68900
rect 206880 68880 207120 68900
rect 207380 68880 207620 68900
rect 207880 68880 208000 68900
rect 196000 68850 196100 68880
rect 196000 68650 196020 68850
rect 196090 68650 196100 68850
rect 196000 68620 196100 68650
rect 196400 68850 196600 68880
rect 196400 68650 196410 68850
rect 196480 68650 196520 68850
rect 196590 68650 196600 68850
rect 196400 68620 196600 68650
rect 196900 68850 197100 68880
rect 196900 68650 196910 68850
rect 196980 68650 197020 68850
rect 197090 68650 197100 68850
rect 196900 68620 197100 68650
rect 197400 68850 197600 68880
rect 197400 68650 197410 68850
rect 197480 68650 197520 68850
rect 197590 68650 197600 68850
rect 197400 68620 197600 68650
rect 197900 68850 198100 68880
rect 197900 68650 197910 68850
rect 197980 68650 198020 68850
rect 198090 68650 198100 68850
rect 197900 68620 198100 68650
rect 198400 68850 198600 68880
rect 198400 68650 198410 68850
rect 198480 68650 198520 68850
rect 198590 68650 198600 68850
rect 198400 68620 198600 68650
rect 198900 68850 199100 68880
rect 198900 68650 198910 68850
rect 198980 68650 199020 68850
rect 199090 68650 199100 68850
rect 198900 68620 199100 68650
rect 199400 68850 199600 68880
rect 199400 68650 199410 68850
rect 199480 68650 199520 68850
rect 199590 68650 199600 68850
rect 199400 68620 199600 68650
rect 199900 68850 200100 68880
rect 199900 68650 199910 68850
rect 199980 68650 200020 68850
rect 200090 68650 200100 68850
rect 199900 68620 200100 68650
rect 200400 68850 200600 68880
rect 200400 68650 200410 68850
rect 200480 68650 200520 68850
rect 200590 68650 200600 68850
rect 200400 68620 200600 68650
rect 200900 68850 201100 68880
rect 200900 68650 200910 68850
rect 200980 68650 201020 68850
rect 201090 68650 201100 68850
rect 200900 68620 201100 68650
rect 201400 68850 201600 68880
rect 201400 68650 201410 68850
rect 201480 68650 201520 68850
rect 201590 68650 201600 68850
rect 201400 68620 201600 68650
rect 201900 68850 202100 68880
rect 201900 68650 201910 68850
rect 201980 68650 202020 68850
rect 202090 68650 202100 68850
rect 201900 68620 202100 68650
rect 202400 68850 202600 68880
rect 202400 68650 202410 68850
rect 202480 68650 202520 68850
rect 202590 68650 202600 68850
rect 202400 68620 202600 68650
rect 202900 68850 203100 68880
rect 202900 68650 202910 68850
rect 202980 68650 203020 68850
rect 203090 68650 203100 68850
rect 202900 68620 203100 68650
rect 203400 68850 203600 68880
rect 203400 68650 203410 68850
rect 203480 68650 203520 68850
rect 203590 68650 203600 68850
rect 203400 68620 203600 68650
rect 203900 68850 204100 68880
rect 203900 68650 203910 68850
rect 203980 68650 204020 68850
rect 204090 68650 204100 68850
rect 203900 68620 204100 68650
rect 204400 68850 204600 68880
rect 204400 68650 204410 68850
rect 204480 68650 204520 68850
rect 204590 68650 204600 68850
rect 204400 68620 204600 68650
rect 204900 68850 205100 68880
rect 204900 68650 204910 68850
rect 204980 68650 205020 68850
rect 205090 68650 205100 68850
rect 204900 68620 205100 68650
rect 205400 68850 205600 68880
rect 205400 68650 205410 68850
rect 205480 68650 205520 68850
rect 205590 68650 205600 68850
rect 205400 68620 205600 68650
rect 205900 68850 206100 68880
rect 205900 68650 205910 68850
rect 205980 68650 206020 68850
rect 206090 68650 206100 68850
rect 205900 68620 206100 68650
rect 206400 68850 206600 68880
rect 206400 68650 206410 68850
rect 206480 68650 206520 68850
rect 206590 68650 206600 68850
rect 206400 68620 206600 68650
rect 206900 68850 207100 68880
rect 206900 68650 206910 68850
rect 206980 68650 207020 68850
rect 207090 68650 207100 68850
rect 206900 68620 207100 68650
rect 207400 68850 207600 68880
rect 207400 68650 207410 68850
rect 207480 68650 207520 68850
rect 207590 68650 207600 68850
rect 207400 68620 207600 68650
rect 207900 68850 208000 68880
rect 207900 68650 207910 68850
rect 207980 68650 208000 68850
rect 207900 68620 208000 68650
rect 196000 68600 196120 68620
rect 196380 68600 196620 68620
rect 196880 68600 197120 68620
rect 197380 68600 197620 68620
rect 197880 68600 198120 68620
rect 198380 68600 198620 68620
rect 198880 68600 199120 68620
rect 199380 68600 199620 68620
rect 199880 68600 200120 68620
rect 200380 68600 200620 68620
rect 200880 68600 201120 68620
rect 201380 68600 201620 68620
rect 201880 68600 202120 68620
rect 202380 68600 202620 68620
rect 202880 68600 203120 68620
rect 203380 68600 203620 68620
rect 203880 68600 204120 68620
rect 204380 68600 204620 68620
rect 204880 68600 205120 68620
rect 205380 68600 205620 68620
rect 205880 68600 206120 68620
rect 206380 68600 206620 68620
rect 206880 68600 207120 68620
rect 207380 68600 207620 68620
rect 207880 68600 208000 68620
rect 196000 68590 208000 68600
rect 196000 68520 196150 68590
rect 196350 68520 196650 68590
rect 196850 68520 197150 68590
rect 197350 68520 197650 68590
rect 197850 68520 198150 68590
rect 198350 68520 198650 68590
rect 198850 68520 199150 68590
rect 199350 68520 199650 68590
rect 199850 68520 200150 68590
rect 200350 68520 200650 68590
rect 200850 68520 201150 68590
rect 201350 68520 201650 68590
rect 201850 68520 202150 68590
rect 202350 68520 202650 68590
rect 202850 68520 203150 68590
rect 203350 68520 203650 68590
rect 203850 68520 204150 68590
rect 204350 68520 204650 68590
rect 204850 68520 205150 68590
rect 205350 68520 205650 68590
rect 205850 68520 206150 68590
rect 206350 68520 206650 68590
rect 206850 68520 207150 68590
rect 207350 68520 207650 68590
rect 207850 68520 208000 68590
rect 196000 68480 208000 68520
rect 196000 68410 196150 68480
rect 196350 68410 196650 68480
rect 196850 68410 197150 68480
rect 197350 68410 197650 68480
rect 197850 68410 198150 68480
rect 198350 68410 198650 68480
rect 198850 68410 199150 68480
rect 199350 68410 199650 68480
rect 199850 68410 200150 68480
rect 200350 68410 200650 68480
rect 200850 68410 201150 68480
rect 201350 68410 201650 68480
rect 201850 68410 202150 68480
rect 202350 68410 202650 68480
rect 202850 68410 203150 68480
rect 203350 68410 203650 68480
rect 203850 68410 204150 68480
rect 204350 68410 204650 68480
rect 204850 68410 205150 68480
rect 205350 68410 205650 68480
rect 205850 68410 206150 68480
rect 206350 68410 206650 68480
rect 206850 68410 207150 68480
rect 207350 68410 207650 68480
rect 207850 68410 208000 68480
rect 196000 68400 208000 68410
rect 196000 68380 196120 68400
rect 196380 68380 196620 68400
rect 196880 68380 197120 68400
rect 197380 68380 197620 68400
rect 197880 68380 198120 68400
rect 198380 68380 198620 68400
rect 198880 68380 199120 68400
rect 199380 68380 199620 68400
rect 199880 68380 200120 68400
rect 200380 68380 200620 68400
rect 200880 68380 201120 68400
rect 201380 68380 201620 68400
rect 201880 68380 202120 68400
rect 202380 68380 202620 68400
rect 202880 68380 203120 68400
rect 203380 68380 203620 68400
rect 203880 68380 204120 68400
rect 204380 68380 204620 68400
rect 204880 68380 205120 68400
rect 205380 68380 205620 68400
rect 205880 68380 206120 68400
rect 206380 68380 206620 68400
rect 206880 68380 207120 68400
rect 207380 68380 207620 68400
rect 207880 68380 208000 68400
rect 196000 68350 196100 68380
rect 196000 68150 196020 68350
rect 196090 68150 196100 68350
rect 196000 68120 196100 68150
rect 196400 68350 196600 68380
rect 196400 68150 196410 68350
rect 196480 68150 196520 68350
rect 196590 68150 196600 68350
rect 196400 68120 196600 68150
rect 196900 68350 197100 68380
rect 196900 68150 196910 68350
rect 196980 68150 197020 68350
rect 197090 68150 197100 68350
rect 196900 68120 197100 68150
rect 197400 68350 197600 68380
rect 197400 68150 197410 68350
rect 197480 68150 197520 68350
rect 197590 68150 197600 68350
rect 197400 68120 197600 68150
rect 197900 68350 198100 68380
rect 197900 68150 197910 68350
rect 197980 68150 198020 68350
rect 198090 68150 198100 68350
rect 197900 68120 198100 68150
rect 198400 68350 198600 68380
rect 198400 68150 198410 68350
rect 198480 68150 198520 68350
rect 198590 68150 198600 68350
rect 198400 68120 198600 68150
rect 198900 68350 199100 68380
rect 198900 68150 198910 68350
rect 198980 68150 199020 68350
rect 199090 68150 199100 68350
rect 198900 68120 199100 68150
rect 199400 68350 199600 68380
rect 199400 68150 199410 68350
rect 199480 68150 199520 68350
rect 199590 68150 199600 68350
rect 199400 68120 199600 68150
rect 199900 68350 200100 68380
rect 199900 68150 199910 68350
rect 199980 68150 200020 68350
rect 200090 68150 200100 68350
rect 199900 68120 200100 68150
rect 200400 68350 200600 68380
rect 200400 68150 200410 68350
rect 200480 68150 200520 68350
rect 200590 68150 200600 68350
rect 200400 68120 200600 68150
rect 200900 68350 201100 68380
rect 200900 68150 200910 68350
rect 200980 68150 201020 68350
rect 201090 68150 201100 68350
rect 200900 68120 201100 68150
rect 201400 68350 201600 68380
rect 201400 68150 201410 68350
rect 201480 68150 201520 68350
rect 201590 68150 201600 68350
rect 201400 68120 201600 68150
rect 201900 68350 202100 68380
rect 201900 68150 201910 68350
rect 201980 68150 202020 68350
rect 202090 68150 202100 68350
rect 201900 68120 202100 68150
rect 202400 68350 202600 68380
rect 202400 68150 202410 68350
rect 202480 68150 202520 68350
rect 202590 68150 202600 68350
rect 202400 68120 202600 68150
rect 202900 68350 203100 68380
rect 202900 68150 202910 68350
rect 202980 68150 203020 68350
rect 203090 68150 203100 68350
rect 202900 68120 203100 68150
rect 203400 68350 203600 68380
rect 203400 68150 203410 68350
rect 203480 68150 203520 68350
rect 203590 68150 203600 68350
rect 203400 68120 203600 68150
rect 203900 68350 204100 68380
rect 203900 68150 203910 68350
rect 203980 68150 204020 68350
rect 204090 68150 204100 68350
rect 203900 68120 204100 68150
rect 204400 68350 204600 68380
rect 204400 68150 204410 68350
rect 204480 68150 204520 68350
rect 204590 68150 204600 68350
rect 204400 68120 204600 68150
rect 204900 68350 205100 68380
rect 204900 68150 204910 68350
rect 204980 68150 205020 68350
rect 205090 68150 205100 68350
rect 204900 68120 205100 68150
rect 205400 68350 205600 68380
rect 205400 68150 205410 68350
rect 205480 68150 205520 68350
rect 205590 68150 205600 68350
rect 205400 68120 205600 68150
rect 205900 68350 206100 68380
rect 205900 68150 205910 68350
rect 205980 68150 206020 68350
rect 206090 68150 206100 68350
rect 205900 68120 206100 68150
rect 206400 68350 206600 68380
rect 206400 68150 206410 68350
rect 206480 68150 206520 68350
rect 206590 68150 206600 68350
rect 206400 68120 206600 68150
rect 206900 68350 207100 68380
rect 206900 68150 206910 68350
rect 206980 68150 207020 68350
rect 207090 68150 207100 68350
rect 206900 68120 207100 68150
rect 207400 68350 207600 68380
rect 207400 68150 207410 68350
rect 207480 68150 207520 68350
rect 207590 68150 207600 68350
rect 207400 68120 207600 68150
rect 207900 68350 208000 68380
rect 207900 68150 207910 68350
rect 207980 68150 208000 68350
rect 207900 68120 208000 68150
rect 196000 68100 196120 68120
rect 196380 68100 196620 68120
rect 196880 68100 197120 68120
rect 197380 68100 197620 68120
rect 197880 68100 198120 68120
rect 198380 68100 198620 68120
rect 198880 68100 199120 68120
rect 199380 68100 199620 68120
rect 199880 68100 200120 68120
rect 200380 68100 200620 68120
rect 200880 68100 201120 68120
rect 201380 68100 201620 68120
rect 201880 68100 202120 68120
rect 202380 68100 202620 68120
rect 202880 68100 203120 68120
rect 203380 68100 203620 68120
rect 203880 68100 204120 68120
rect 204380 68100 204620 68120
rect 204880 68100 205120 68120
rect 205380 68100 205620 68120
rect 205880 68100 206120 68120
rect 206380 68100 206620 68120
rect 206880 68100 207120 68120
rect 207380 68100 207620 68120
rect 207880 68100 208000 68120
rect 196000 68090 208000 68100
rect 196000 68020 196150 68090
rect 196350 68020 196650 68090
rect 196850 68020 197150 68090
rect 197350 68020 197650 68090
rect 197850 68020 198150 68090
rect 198350 68020 198650 68090
rect 198850 68020 199150 68090
rect 199350 68020 199650 68090
rect 199850 68020 200150 68090
rect 200350 68020 200650 68090
rect 200850 68020 201150 68090
rect 201350 68020 201650 68090
rect 201850 68020 202150 68090
rect 202350 68020 202650 68090
rect 202850 68020 203150 68090
rect 203350 68020 203650 68090
rect 203850 68020 204150 68090
rect 204350 68020 204650 68090
rect 204850 68020 205150 68090
rect 205350 68020 205650 68090
rect 205850 68020 206150 68090
rect 206350 68020 206650 68090
rect 206850 68020 207150 68090
rect 207350 68020 207650 68090
rect 207850 68020 208000 68090
rect 130000 67900 132000 68000
rect 130000 67880 130120 67900
rect 130380 67880 130620 67900
rect 130880 67880 131120 67900
rect 131380 67880 131620 67900
rect 131880 67880 132000 67900
rect 130000 67620 130100 67880
rect 130400 67620 130600 67880
rect 130900 67620 131100 67880
rect 131400 67620 131600 67880
rect 131900 67620 132000 67880
rect 130000 67600 130120 67620
rect 130380 67600 130620 67620
rect 130880 67600 131120 67620
rect 131380 67600 131620 67620
rect 131880 67600 132000 67620
rect 130000 67400 132000 67600
rect 130000 67380 130120 67400
rect 130380 67380 130620 67400
rect 130880 67380 131120 67400
rect 131380 67380 131620 67400
rect 131880 67380 132000 67400
rect 130000 67120 130100 67380
rect 130400 67120 130600 67380
rect 130900 67120 131100 67380
rect 131400 67120 131600 67380
rect 131900 67120 132000 67380
rect 130000 67100 130120 67120
rect 130380 67100 130620 67120
rect 130880 67100 131120 67120
rect 131380 67100 131620 67120
rect 131880 67100 132000 67120
rect 130000 66900 132000 67100
rect 130000 66880 130120 66900
rect 130380 66880 130620 66900
rect 130880 66880 131120 66900
rect 131380 66880 131620 66900
rect 131880 66880 132000 66900
rect 130000 66620 130100 66880
rect 130400 66620 130600 66880
rect 130900 66620 131100 66880
rect 131400 66620 131600 66880
rect 131900 66620 132000 66880
rect 130000 66600 130120 66620
rect 130380 66600 130620 66620
rect 130880 66600 131120 66620
rect 131380 66600 131620 66620
rect 131880 66600 132000 66620
rect 130000 66400 132000 66600
rect 130000 66380 130120 66400
rect 130380 66380 130620 66400
rect 130880 66380 131120 66400
rect 131380 66380 131620 66400
rect 131880 66380 132000 66400
rect 130000 66120 130100 66380
rect 130400 66120 130600 66380
rect 130900 66120 131100 66380
rect 131400 66120 131600 66380
rect 131900 66120 132000 66380
rect 130000 66100 130120 66120
rect 130380 66100 130620 66120
rect 130880 66100 131120 66120
rect 131380 66100 131620 66120
rect 131880 66100 132000 66120
rect 130000 65900 132000 66100
rect 196000 67980 208000 68020
rect 196000 67910 196150 67980
rect 196350 67910 196650 67980
rect 196850 67910 197150 67980
rect 197350 67910 197650 67980
rect 197850 67910 198150 67980
rect 198350 67910 198650 67980
rect 198850 67910 199150 67980
rect 199350 67910 199650 67980
rect 199850 67910 200150 67980
rect 200350 67910 200650 67980
rect 200850 67910 201150 67980
rect 201350 67910 201650 67980
rect 201850 67910 202150 67980
rect 202350 67910 202650 67980
rect 202850 67910 203150 67980
rect 203350 67910 203650 67980
rect 203850 67910 204150 67980
rect 204350 67910 204650 67980
rect 204850 67910 205150 67980
rect 205350 67910 205650 67980
rect 205850 67910 206150 67980
rect 206350 67910 206650 67980
rect 206850 67910 207150 67980
rect 207350 67910 207650 67980
rect 207850 67910 208000 67980
rect 196000 67900 208000 67910
rect 196000 67880 196120 67900
rect 196380 67880 196620 67900
rect 196880 67880 197120 67900
rect 197380 67880 197620 67900
rect 197880 67880 198120 67900
rect 198380 67880 198620 67900
rect 198880 67880 199120 67900
rect 199380 67880 199620 67900
rect 199880 67880 200120 67900
rect 200380 67880 200620 67900
rect 200880 67880 201120 67900
rect 201380 67880 201620 67900
rect 201880 67880 202120 67900
rect 202380 67880 202620 67900
rect 202880 67880 203120 67900
rect 203380 67880 203620 67900
rect 203880 67880 204120 67900
rect 204380 67880 204620 67900
rect 204880 67880 205120 67900
rect 205380 67880 205620 67900
rect 205880 67880 206120 67900
rect 206380 67880 206620 67900
rect 206880 67880 207120 67900
rect 207380 67880 207620 67900
rect 207880 67880 208000 67900
rect 196000 67850 196100 67880
rect 196000 67650 196020 67850
rect 196090 67650 196100 67850
rect 196000 67620 196100 67650
rect 196400 67850 196600 67880
rect 196400 67650 196410 67850
rect 196480 67650 196520 67850
rect 196590 67650 196600 67850
rect 196400 67620 196600 67650
rect 196900 67850 197100 67880
rect 196900 67650 196910 67850
rect 196980 67650 197020 67850
rect 197090 67650 197100 67850
rect 196900 67620 197100 67650
rect 197400 67850 197600 67880
rect 197400 67650 197410 67850
rect 197480 67650 197520 67850
rect 197590 67650 197600 67850
rect 197400 67620 197600 67650
rect 197900 67850 198100 67880
rect 197900 67650 197910 67850
rect 197980 67650 198020 67850
rect 198090 67650 198100 67850
rect 197900 67620 198100 67650
rect 198400 67850 198600 67880
rect 198400 67650 198410 67850
rect 198480 67650 198520 67850
rect 198590 67650 198600 67850
rect 198400 67620 198600 67650
rect 198900 67850 199100 67880
rect 198900 67650 198910 67850
rect 198980 67650 199020 67850
rect 199090 67650 199100 67850
rect 198900 67620 199100 67650
rect 199400 67850 199600 67880
rect 199400 67650 199410 67850
rect 199480 67650 199520 67850
rect 199590 67650 199600 67850
rect 199400 67620 199600 67650
rect 199900 67850 200100 67880
rect 199900 67650 199910 67850
rect 199980 67650 200020 67850
rect 200090 67650 200100 67850
rect 199900 67620 200100 67650
rect 200400 67850 200600 67880
rect 200400 67650 200410 67850
rect 200480 67650 200520 67850
rect 200590 67650 200600 67850
rect 200400 67620 200600 67650
rect 200900 67850 201100 67880
rect 200900 67650 200910 67850
rect 200980 67650 201020 67850
rect 201090 67650 201100 67850
rect 200900 67620 201100 67650
rect 201400 67850 201600 67880
rect 201400 67650 201410 67850
rect 201480 67650 201520 67850
rect 201590 67650 201600 67850
rect 201400 67620 201600 67650
rect 201900 67850 202100 67880
rect 201900 67650 201910 67850
rect 201980 67650 202020 67850
rect 202090 67650 202100 67850
rect 201900 67620 202100 67650
rect 202400 67850 202600 67880
rect 202400 67650 202410 67850
rect 202480 67650 202520 67850
rect 202590 67650 202600 67850
rect 202400 67620 202600 67650
rect 202900 67850 203100 67880
rect 202900 67650 202910 67850
rect 202980 67650 203020 67850
rect 203090 67650 203100 67850
rect 202900 67620 203100 67650
rect 203400 67850 203600 67880
rect 203400 67650 203410 67850
rect 203480 67650 203520 67850
rect 203590 67650 203600 67850
rect 203400 67620 203600 67650
rect 203900 67850 204100 67880
rect 203900 67650 203910 67850
rect 203980 67650 204020 67850
rect 204090 67650 204100 67850
rect 203900 67620 204100 67650
rect 204400 67850 204600 67880
rect 204400 67650 204410 67850
rect 204480 67650 204520 67850
rect 204590 67650 204600 67850
rect 204400 67620 204600 67650
rect 204900 67850 205100 67880
rect 204900 67650 204910 67850
rect 204980 67650 205020 67850
rect 205090 67650 205100 67850
rect 204900 67620 205100 67650
rect 205400 67850 205600 67880
rect 205400 67650 205410 67850
rect 205480 67650 205520 67850
rect 205590 67650 205600 67850
rect 205400 67620 205600 67650
rect 205900 67850 206100 67880
rect 205900 67650 205910 67850
rect 205980 67650 206020 67850
rect 206090 67650 206100 67850
rect 205900 67620 206100 67650
rect 206400 67850 206600 67880
rect 206400 67650 206410 67850
rect 206480 67650 206520 67850
rect 206590 67650 206600 67850
rect 206400 67620 206600 67650
rect 206900 67850 207100 67880
rect 206900 67650 206910 67850
rect 206980 67650 207020 67850
rect 207090 67650 207100 67850
rect 206900 67620 207100 67650
rect 207400 67850 207600 67880
rect 207400 67650 207410 67850
rect 207480 67650 207520 67850
rect 207590 67650 207600 67850
rect 207400 67620 207600 67650
rect 207900 67850 208000 67880
rect 207900 67650 207910 67850
rect 207980 67650 208000 67850
rect 207900 67620 208000 67650
rect 196000 67600 196120 67620
rect 196380 67600 196620 67620
rect 196880 67600 197120 67620
rect 197380 67600 197620 67620
rect 197880 67600 198120 67620
rect 198380 67600 198620 67620
rect 198880 67600 199120 67620
rect 199380 67600 199620 67620
rect 199880 67600 200120 67620
rect 200380 67600 200620 67620
rect 200880 67600 201120 67620
rect 201380 67600 201620 67620
rect 201880 67600 202120 67620
rect 202380 67600 202620 67620
rect 202880 67600 203120 67620
rect 203380 67600 203620 67620
rect 203880 67600 204120 67620
rect 204380 67600 204620 67620
rect 204880 67600 205120 67620
rect 205380 67600 205620 67620
rect 205880 67600 206120 67620
rect 206380 67600 206620 67620
rect 206880 67600 207120 67620
rect 207380 67600 207620 67620
rect 207880 67600 208000 67620
rect 196000 67590 208000 67600
rect 196000 67520 196150 67590
rect 196350 67520 196650 67590
rect 196850 67520 197150 67590
rect 197350 67520 197650 67590
rect 197850 67520 198150 67590
rect 198350 67520 198650 67590
rect 198850 67520 199150 67590
rect 199350 67520 199650 67590
rect 199850 67520 200150 67590
rect 200350 67520 200650 67590
rect 200850 67520 201150 67590
rect 201350 67520 201650 67590
rect 201850 67520 202150 67590
rect 202350 67520 202650 67590
rect 202850 67520 203150 67590
rect 203350 67520 203650 67590
rect 203850 67520 204150 67590
rect 204350 67520 204650 67590
rect 204850 67520 205150 67590
rect 205350 67520 205650 67590
rect 205850 67520 206150 67590
rect 206350 67520 206650 67590
rect 206850 67520 207150 67590
rect 207350 67520 207650 67590
rect 207850 67520 208000 67590
rect 196000 67480 208000 67520
rect 196000 67410 196150 67480
rect 196350 67410 196650 67480
rect 196850 67410 197150 67480
rect 197350 67410 197650 67480
rect 197850 67410 198150 67480
rect 198350 67410 198650 67480
rect 198850 67410 199150 67480
rect 199350 67410 199650 67480
rect 199850 67410 200150 67480
rect 200350 67410 200650 67480
rect 200850 67410 201150 67480
rect 201350 67410 201650 67480
rect 201850 67410 202150 67480
rect 202350 67410 202650 67480
rect 202850 67410 203150 67480
rect 203350 67410 203650 67480
rect 203850 67410 204150 67480
rect 204350 67410 204650 67480
rect 204850 67410 205150 67480
rect 205350 67410 205650 67480
rect 205850 67410 206150 67480
rect 206350 67410 206650 67480
rect 206850 67410 207150 67480
rect 207350 67410 207650 67480
rect 207850 67410 208000 67480
rect 196000 67400 208000 67410
rect 196000 67380 196120 67400
rect 196380 67380 196620 67400
rect 196880 67380 197120 67400
rect 197380 67380 197620 67400
rect 197880 67380 198120 67400
rect 198380 67380 198620 67400
rect 198880 67380 199120 67400
rect 199380 67380 199620 67400
rect 199880 67380 200120 67400
rect 200380 67380 200620 67400
rect 200880 67380 201120 67400
rect 201380 67380 201620 67400
rect 201880 67380 202120 67400
rect 202380 67380 202620 67400
rect 202880 67380 203120 67400
rect 203380 67380 203620 67400
rect 203880 67380 204120 67400
rect 204380 67380 204620 67400
rect 204880 67380 205120 67400
rect 205380 67380 205620 67400
rect 205880 67380 206120 67400
rect 206380 67380 206620 67400
rect 206880 67380 207120 67400
rect 207380 67380 207620 67400
rect 207880 67380 208000 67400
rect 196000 67350 196100 67380
rect 196000 67150 196020 67350
rect 196090 67150 196100 67350
rect 196000 67120 196100 67150
rect 196400 67350 196600 67380
rect 196400 67150 196410 67350
rect 196480 67150 196520 67350
rect 196590 67150 196600 67350
rect 196400 67120 196600 67150
rect 196900 67350 197100 67380
rect 196900 67150 196910 67350
rect 196980 67150 197020 67350
rect 197090 67150 197100 67350
rect 196900 67120 197100 67150
rect 197400 67350 197600 67380
rect 197400 67150 197410 67350
rect 197480 67150 197520 67350
rect 197590 67150 197600 67350
rect 197400 67120 197600 67150
rect 197900 67350 198100 67380
rect 197900 67150 197910 67350
rect 197980 67150 198020 67350
rect 198090 67150 198100 67350
rect 197900 67120 198100 67150
rect 198400 67350 198600 67380
rect 198400 67150 198410 67350
rect 198480 67150 198520 67350
rect 198590 67150 198600 67350
rect 198400 67120 198600 67150
rect 198900 67350 199100 67380
rect 198900 67150 198910 67350
rect 198980 67150 199020 67350
rect 199090 67150 199100 67350
rect 198900 67120 199100 67150
rect 199400 67350 199600 67380
rect 199400 67150 199410 67350
rect 199480 67150 199520 67350
rect 199590 67150 199600 67350
rect 199400 67120 199600 67150
rect 199900 67350 200100 67380
rect 199900 67150 199910 67350
rect 199980 67150 200020 67350
rect 200090 67150 200100 67350
rect 199900 67120 200100 67150
rect 200400 67350 200600 67380
rect 200400 67150 200410 67350
rect 200480 67150 200520 67350
rect 200590 67150 200600 67350
rect 200400 67120 200600 67150
rect 200900 67350 201100 67380
rect 200900 67150 200910 67350
rect 200980 67150 201020 67350
rect 201090 67150 201100 67350
rect 200900 67120 201100 67150
rect 201400 67350 201600 67380
rect 201400 67150 201410 67350
rect 201480 67150 201520 67350
rect 201590 67150 201600 67350
rect 201400 67120 201600 67150
rect 201900 67350 202100 67380
rect 201900 67150 201910 67350
rect 201980 67150 202020 67350
rect 202090 67150 202100 67350
rect 201900 67120 202100 67150
rect 202400 67350 202600 67380
rect 202400 67150 202410 67350
rect 202480 67150 202520 67350
rect 202590 67150 202600 67350
rect 202400 67120 202600 67150
rect 202900 67350 203100 67380
rect 202900 67150 202910 67350
rect 202980 67150 203020 67350
rect 203090 67150 203100 67350
rect 202900 67120 203100 67150
rect 203400 67350 203600 67380
rect 203400 67150 203410 67350
rect 203480 67150 203520 67350
rect 203590 67150 203600 67350
rect 203400 67120 203600 67150
rect 203900 67350 204100 67380
rect 203900 67150 203910 67350
rect 203980 67150 204020 67350
rect 204090 67150 204100 67350
rect 203900 67120 204100 67150
rect 204400 67350 204600 67380
rect 204400 67150 204410 67350
rect 204480 67150 204520 67350
rect 204590 67150 204600 67350
rect 204400 67120 204600 67150
rect 204900 67350 205100 67380
rect 204900 67150 204910 67350
rect 204980 67150 205020 67350
rect 205090 67150 205100 67350
rect 204900 67120 205100 67150
rect 205400 67350 205600 67380
rect 205400 67150 205410 67350
rect 205480 67150 205520 67350
rect 205590 67150 205600 67350
rect 205400 67120 205600 67150
rect 205900 67350 206100 67380
rect 205900 67150 205910 67350
rect 205980 67150 206020 67350
rect 206090 67150 206100 67350
rect 205900 67120 206100 67150
rect 206400 67350 206600 67380
rect 206400 67150 206410 67350
rect 206480 67150 206520 67350
rect 206590 67150 206600 67350
rect 206400 67120 206600 67150
rect 206900 67350 207100 67380
rect 206900 67150 206910 67350
rect 206980 67150 207020 67350
rect 207090 67150 207100 67350
rect 206900 67120 207100 67150
rect 207400 67350 207600 67380
rect 207400 67150 207410 67350
rect 207480 67150 207520 67350
rect 207590 67150 207600 67350
rect 207400 67120 207600 67150
rect 207900 67350 208000 67380
rect 207900 67150 207910 67350
rect 207980 67150 208000 67350
rect 207900 67120 208000 67150
rect 196000 67100 196120 67120
rect 196380 67100 196620 67120
rect 196880 67100 197120 67120
rect 197380 67100 197620 67120
rect 197880 67100 198120 67120
rect 198380 67100 198620 67120
rect 198880 67100 199120 67120
rect 199380 67100 199620 67120
rect 199880 67100 200120 67120
rect 200380 67100 200620 67120
rect 200880 67100 201120 67120
rect 201380 67100 201620 67120
rect 201880 67100 202120 67120
rect 202380 67100 202620 67120
rect 202880 67100 203120 67120
rect 203380 67100 203620 67120
rect 203880 67100 204120 67120
rect 204380 67100 204620 67120
rect 204880 67100 205120 67120
rect 205380 67100 205620 67120
rect 205880 67100 206120 67120
rect 206380 67100 206620 67120
rect 206880 67100 207120 67120
rect 207380 67100 207620 67120
rect 207880 67100 208000 67120
rect 196000 67090 208000 67100
rect 196000 67020 196150 67090
rect 196350 67020 196650 67090
rect 196850 67020 197150 67090
rect 197350 67020 197650 67090
rect 197850 67020 198150 67090
rect 198350 67020 198650 67090
rect 198850 67020 199150 67090
rect 199350 67020 199650 67090
rect 199850 67020 200150 67090
rect 200350 67020 200650 67090
rect 200850 67020 201150 67090
rect 201350 67020 201650 67090
rect 201850 67020 202150 67090
rect 202350 67020 202650 67090
rect 202850 67020 203150 67090
rect 203350 67020 203650 67090
rect 203850 67020 204150 67090
rect 204350 67020 204650 67090
rect 204850 67020 205150 67090
rect 205350 67020 205650 67090
rect 205850 67020 206150 67090
rect 206350 67020 206650 67090
rect 206850 67020 207150 67090
rect 207350 67020 207650 67090
rect 207850 67020 208000 67090
rect 196000 66980 208000 67020
rect 196000 66910 196150 66980
rect 196350 66910 196650 66980
rect 196850 66910 197150 66980
rect 197350 66910 197650 66980
rect 197850 66910 198150 66980
rect 198350 66910 198650 66980
rect 198850 66910 199150 66980
rect 199350 66910 199650 66980
rect 199850 66910 200150 66980
rect 200350 66910 200650 66980
rect 200850 66910 201150 66980
rect 201350 66910 201650 66980
rect 201850 66910 202150 66980
rect 202350 66910 202650 66980
rect 202850 66910 203150 66980
rect 203350 66910 203650 66980
rect 203850 66910 204150 66980
rect 204350 66910 204650 66980
rect 204850 66910 205150 66980
rect 205350 66910 205650 66980
rect 205850 66910 206150 66980
rect 206350 66910 206650 66980
rect 206850 66910 207150 66980
rect 207350 66910 207650 66980
rect 207850 66910 208000 66980
rect 196000 66900 208000 66910
rect 196000 66880 196120 66900
rect 196380 66880 196620 66900
rect 196880 66880 197120 66900
rect 197380 66880 197620 66900
rect 197880 66880 198120 66900
rect 198380 66880 198620 66900
rect 198880 66880 199120 66900
rect 199380 66880 199620 66900
rect 199880 66880 200120 66900
rect 200380 66880 200620 66900
rect 200880 66880 201120 66900
rect 201380 66880 201620 66900
rect 201880 66880 202120 66900
rect 202380 66880 202620 66900
rect 202880 66880 203120 66900
rect 203380 66880 203620 66900
rect 203880 66880 204120 66900
rect 204380 66880 204620 66900
rect 204880 66880 205120 66900
rect 205380 66880 205620 66900
rect 205880 66880 206120 66900
rect 206380 66880 206620 66900
rect 206880 66880 207120 66900
rect 207380 66880 207620 66900
rect 207880 66880 208000 66900
rect 196000 66850 196100 66880
rect 196000 66650 196020 66850
rect 196090 66650 196100 66850
rect 196000 66620 196100 66650
rect 196400 66850 196600 66880
rect 196400 66650 196410 66850
rect 196480 66650 196520 66850
rect 196590 66650 196600 66850
rect 196400 66620 196600 66650
rect 196900 66850 197100 66880
rect 196900 66650 196910 66850
rect 196980 66650 197020 66850
rect 197090 66650 197100 66850
rect 196900 66620 197100 66650
rect 197400 66850 197600 66880
rect 197400 66650 197410 66850
rect 197480 66650 197520 66850
rect 197590 66650 197600 66850
rect 197400 66620 197600 66650
rect 197900 66850 198100 66880
rect 197900 66650 197910 66850
rect 197980 66650 198020 66850
rect 198090 66650 198100 66850
rect 197900 66620 198100 66650
rect 198400 66850 198600 66880
rect 198400 66650 198410 66850
rect 198480 66650 198520 66850
rect 198590 66650 198600 66850
rect 198400 66620 198600 66650
rect 198900 66850 199100 66880
rect 198900 66650 198910 66850
rect 198980 66650 199020 66850
rect 199090 66650 199100 66850
rect 198900 66620 199100 66650
rect 199400 66850 199600 66880
rect 199400 66650 199410 66850
rect 199480 66650 199520 66850
rect 199590 66650 199600 66850
rect 199400 66620 199600 66650
rect 199900 66850 200100 66880
rect 199900 66650 199910 66850
rect 199980 66650 200020 66850
rect 200090 66650 200100 66850
rect 199900 66620 200100 66650
rect 200400 66850 200600 66880
rect 200400 66650 200410 66850
rect 200480 66650 200520 66850
rect 200590 66650 200600 66850
rect 200400 66620 200600 66650
rect 200900 66850 201100 66880
rect 200900 66650 200910 66850
rect 200980 66650 201020 66850
rect 201090 66650 201100 66850
rect 200900 66620 201100 66650
rect 201400 66850 201600 66880
rect 201400 66650 201410 66850
rect 201480 66650 201520 66850
rect 201590 66650 201600 66850
rect 201400 66620 201600 66650
rect 201900 66850 202100 66880
rect 201900 66650 201910 66850
rect 201980 66650 202020 66850
rect 202090 66650 202100 66850
rect 201900 66620 202100 66650
rect 202400 66850 202600 66880
rect 202400 66650 202410 66850
rect 202480 66650 202520 66850
rect 202590 66650 202600 66850
rect 202400 66620 202600 66650
rect 202900 66850 203100 66880
rect 202900 66650 202910 66850
rect 202980 66650 203020 66850
rect 203090 66650 203100 66850
rect 202900 66620 203100 66650
rect 203400 66850 203600 66880
rect 203400 66650 203410 66850
rect 203480 66650 203520 66850
rect 203590 66650 203600 66850
rect 203400 66620 203600 66650
rect 203900 66850 204100 66880
rect 203900 66650 203910 66850
rect 203980 66650 204020 66850
rect 204090 66650 204100 66850
rect 203900 66620 204100 66650
rect 204400 66850 204600 66880
rect 204400 66650 204410 66850
rect 204480 66650 204520 66850
rect 204590 66650 204600 66850
rect 204400 66620 204600 66650
rect 204900 66850 205100 66880
rect 204900 66650 204910 66850
rect 204980 66650 205020 66850
rect 205090 66650 205100 66850
rect 204900 66620 205100 66650
rect 205400 66850 205600 66880
rect 205400 66650 205410 66850
rect 205480 66650 205520 66850
rect 205590 66650 205600 66850
rect 205400 66620 205600 66650
rect 205900 66850 206100 66880
rect 205900 66650 205910 66850
rect 205980 66650 206020 66850
rect 206090 66650 206100 66850
rect 205900 66620 206100 66650
rect 206400 66850 206600 66880
rect 206400 66650 206410 66850
rect 206480 66650 206520 66850
rect 206590 66650 206600 66850
rect 206400 66620 206600 66650
rect 206900 66850 207100 66880
rect 206900 66650 206910 66850
rect 206980 66650 207020 66850
rect 207090 66650 207100 66850
rect 206900 66620 207100 66650
rect 207400 66850 207600 66880
rect 207400 66650 207410 66850
rect 207480 66650 207520 66850
rect 207590 66650 207600 66850
rect 207400 66620 207600 66650
rect 207900 66850 208000 66880
rect 207900 66650 207910 66850
rect 207980 66650 208000 66850
rect 207900 66620 208000 66650
rect 196000 66600 196120 66620
rect 196380 66600 196620 66620
rect 196880 66600 197120 66620
rect 197380 66600 197620 66620
rect 197880 66600 198120 66620
rect 198380 66600 198620 66620
rect 198880 66600 199120 66620
rect 199380 66600 199620 66620
rect 199880 66600 200120 66620
rect 200380 66600 200620 66620
rect 200880 66600 201120 66620
rect 201380 66600 201620 66620
rect 201880 66600 202120 66620
rect 202380 66600 202620 66620
rect 202880 66600 203120 66620
rect 203380 66600 203620 66620
rect 203880 66600 204120 66620
rect 204380 66600 204620 66620
rect 204880 66600 205120 66620
rect 205380 66600 205620 66620
rect 205880 66600 206120 66620
rect 206380 66600 206620 66620
rect 206880 66600 207120 66620
rect 207380 66600 207620 66620
rect 207880 66600 208000 66620
rect 196000 66590 208000 66600
rect 196000 66520 196150 66590
rect 196350 66520 196650 66590
rect 196850 66520 197150 66590
rect 197350 66520 197650 66590
rect 197850 66520 198150 66590
rect 198350 66520 198650 66590
rect 198850 66520 199150 66590
rect 199350 66520 199650 66590
rect 199850 66520 200150 66590
rect 200350 66520 200650 66590
rect 200850 66520 201150 66590
rect 201350 66520 201650 66590
rect 201850 66520 202150 66590
rect 202350 66520 202650 66590
rect 202850 66520 203150 66590
rect 203350 66520 203650 66590
rect 203850 66520 204150 66590
rect 204350 66520 204650 66590
rect 204850 66520 205150 66590
rect 205350 66520 205650 66590
rect 205850 66520 206150 66590
rect 206350 66520 206650 66590
rect 206850 66520 207150 66590
rect 207350 66520 207650 66590
rect 207850 66520 208000 66590
rect 196000 66480 208000 66520
rect 196000 66410 196150 66480
rect 196350 66410 196650 66480
rect 196850 66410 197150 66480
rect 197350 66410 197650 66480
rect 197850 66410 198150 66480
rect 198350 66410 198650 66480
rect 198850 66410 199150 66480
rect 199350 66410 199650 66480
rect 199850 66410 200150 66480
rect 200350 66410 200650 66480
rect 200850 66410 201150 66480
rect 201350 66410 201650 66480
rect 201850 66410 202150 66480
rect 202350 66410 202650 66480
rect 202850 66410 203150 66480
rect 203350 66410 203650 66480
rect 203850 66410 204150 66480
rect 204350 66410 204650 66480
rect 204850 66410 205150 66480
rect 205350 66410 205650 66480
rect 205850 66410 206150 66480
rect 206350 66410 206650 66480
rect 206850 66410 207150 66480
rect 207350 66410 207650 66480
rect 207850 66410 208000 66480
rect 196000 66400 208000 66410
rect 196000 66380 196120 66400
rect 196380 66380 196620 66400
rect 196880 66380 197120 66400
rect 197380 66380 197620 66400
rect 197880 66380 198120 66400
rect 198380 66380 198620 66400
rect 198880 66380 199120 66400
rect 199380 66380 199620 66400
rect 199880 66380 200120 66400
rect 200380 66380 200620 66400
rect 200880 66380 201120 66400
rect 201380 66380 201620 66400
rect 201880 66380 202120 66400
rect 202380 66380 202620 66400
rect 202880 66380 203120 66400
rect 203380 66380 203620 66400
rect 203880 66380 204120 66400
rect 204380 66380 204620 66400
rect 204880 66380 205120 66400
rect 205380 66380 205620 66400
rect 205880 66380 206120 66400
rect 206380 66380 206620 66400
rect 206880 66380 207120 66400
rect 207380 66380 207620 66400
rect 207880 66380 208000 66400
rect 196000 66350 196100 66380
rect 196000 66150 196020 66350
rect 196090 66150 196100 66350
rect 196000 66120 196100 66150
rect 196400 66350 196600 66380
rect 196400 66150 196410 66350
rect 196480 66150 196520 66350
rect 196590 66150 196600 66350
rect 196400 66120 196600 66150
rect 196900 66350 197100 66380
rect 196900 66150 196910 66350
rect 196980 66150 197020 66350
rect 197090 66150 197100 66350
rect 196900 66120 197100 66150
rect 197400 66350 197600 66380
rect 197400 66150 197410 66350
rect 197480 66150 197520 66350
rect 197590 66150 197600 66350
rect 197400 66120 197600 66150
rect 197900 66350 198100 66380
rect 197900 66150 197910 66350
rect 197980 66150 198020 66350
rect 198090 66150 198100 66350
rect 197900 66120 198100 66150
rect 198400 66350 198600 66380
rect 198400 66150 198410 66350
rect 198480 66150 198520 66350
rect 198590 66150 198600 66350
rect 198400 66120 198600 66150
rect 198900 66350 199100 66380
rect 198900 66150 198910 66350
rect 198980 66150 199020 66350
rect 199090 66150 199100 66350
rect 198900 66120 199100 66150
rect 199400 66350 199600 66380
rect 199400 66150 199410 66350
rect 199480 66150 199520 66350
rect 199590 66150 199600 66350
rect 199400 66120 199600 66150
rect 199900 66350 200100 66380
rect 199900 66150 199910 66350
rect 199980 66150 200020 66350
rect 200090 66150 200100 66350
rect 199900 66120 200100 66150
rect 200400 66350 200600 66380
rect 200400 66150 200410 66350
rect 200480 66150 200520 66350
rect 200590 66150 200600 66350
rect 200400 66120 200600 66150
rect 200900 66350 201100 66380
rect 200900 66150 200910 66350
rect 200980 66150 201020 66350
rect 201090 66150 201100 66350
rect 200900 66120 201100 66150
rect 201400 66350 201600 66380
rect 201400 66150 201410 66350
rect 201480 66150 201520 66350
rect 201590 66150 201600 66350
rect 201400 66120 201600 66150
rect 201900 66350 202100 66380
rect 201900 66150 201910 66350
rect 201980 66150 202020 66350
rect 202090 66150 202100 66350
rect 201900 66120 202100 66150
rect 202400 66350 202600 66380
rect 202400 66150 202410 66350
rect 202480 66150 202520 66350
rect 202590 66150 202600 66350
rect 202400 66120 202600 66150
rect 202900 66350 203100 66380
rect 202900 66150 202910 66350
rect 202980 66150 203020 66350
rect 203090 66150 203100 66350
rect 202900 66120 203100 66150
rect 203400 66350 203600 66380
rect 203400 66150 203410 66350
rect 203480 66150 203520 66350
rect 203590 66150 203600 66350
rect 203400 66120 203600 66150
rect 203900 66350 204100 66380
rect 203900 66150 203910 66350
rect 203980 66150 204020 66350
rect 204090 66150 204100 66350
rect 203900 66120 204100 66150
rect 204400 66350 204600 66380
rect 204400 66150 204410 66350
rect 204480 66150 204520 66350
rect 204590 66150 204600 66350
rect 204400 66120 204600 66150
rect 204900 66350 205100 66380
rect 204900 66150 204910 66350
rect 204980 66150 205020 66350
rect 205090 66150 205100 66350
rect 204900 66120 205100 66150
rect 205400 66350 205600 66380
rect 205400 66150 205410 66350
rect 205480 66150 205520 66350
rect 205590 66150 205600 66350
rect 205400 66120 205600 66150
rect 205900 66350 206100 66380
rect 205900 66150 205910 66350
rect 205980 66150 206020 66350
rect 206090 66150 206100 66350
rect 205900 66120 206100 66150
rect 206400 66350 206600 66380
rect 206400 66150 206410 66350
rect 206480 66150 206520 66350
rect 206590 66150 206600 66350
rect 206400 66120 206600 66150
rect 206900 66350 207100 66380
rect 206900 66150 206910 66350
rect 206980 66150 207020 66350
rect 207090 66150 207100 66350
rect 206900 66120 207100 66150
rect 207400 66350 207600 66380
rect 207400 66150 207410 66350
rect 207480 66150 207520 66350
rect 207590 66150 207600 66350
rect 207400 66120 207600 66150
rect 207900 66350 208000 66380
rect 207900 66150 207910 66350
rect 207980 66150 208000 66350
rect 207900 66120 208000 66150
rect 196000 66100 196120 66120
rect 196380 66100 196620 66120
rect 196880 66100 197120 66120
rect 197380 66100 197620 66120
rect 197880 66100 198120 66120
rect 198380 66100 198620 66120
rect 198880 66100 199120 66120
rect 199380 66100 199620 66120
rect 199880 66100 200120 66120
rect 200380 66100 200620 66120
rect 200880 66100 201120 66120
rect 201380 66100 201620 66120
rect 201880 66100 202120 66120
rect 202380 66100 202620 66120
rect 202880 66100 203120 66120
rect 203380 66100 203620 66120
rect 203880 66100 204120 66120
rect 204380 66100 204620 66120
rect 204880 66100 205120 66120
rect 205380 66100 205620 66120
rect 205880 66100 206120 66120
rect 206380 66100 206620 66120
rect 206880 66100 207120 66120
rect 207380 66100 207620 66120
rect 207880 66100 208000 66120
rect 196000 66090 208000 66100
rect 196000 66020 196150 66090
rect 196350 66020 196650 66090
rect 196850 66020 197150 66090
rect 197350 66020 197650 66090
rect 197850 66020 198150 66090
rect 198350 66020 198650 66090
rect 198850 66020 199150 66090
rect 199350 66020 199650 66090
rect 199850 66020 200150 66090
rect 200350 66020 200650 66090
rect 200850 66020 201150 66090
rect 201350 66020 201650 66090
rect 201850 66020 202150 66090
rect 202350 66020 202650 66090
rect 202850 66020 203150 66090
rect 203350 66020 203650 66090
rect 203850 66020 204150 66090
rect 204350 66020 204650 66090
rect 204850 66020 205150 66090
rect 205350 66020 205650 66090
rect 205850 66020 206150 66090
rect 206350 66020 206650 66090
rect 206850 66020 207150 66090
rect 207350 66020 207650 66090
rect 207850 66020 208000 66090
rect 196000 66000 208000 66020
rect 130000 65880 130120 65900
rect 130380 65880 130620 65900
rect 130880 65880 131120 65900
rect 131380 65880 131620 65900
rect 131880 65880 132000 65900
rect 130000 65620 130100 65880
rect 130400 65620 130600 65880
rect 130900 65620 131100 65880
rect 131400 65620 131600 65880
rect 131900 65620 132000 65880
rect 130000 65600 130120 65620
rect 130380 65600 130620 65620
rect 130880 65600 131120 65620
rect 131380 65600 131620 65620
rect 131880 65600 132000 65620
rect 130000 65400 132000 65600
rect 130000 65380 130120 65400
rect 130380 65380 130620 65400
rect 130880 65380 131120 65400
rect 131380 65380 131620 65400
rect 131880 65380 132000 65400
rect 130000 65120 130100 65380
rect 130400 65120 130600 65380
rect 130900 65120 131100 65380
rect 131400 65120 131600 65380
rect 131900 65120 132000 65380
rect 130000 65100 130120 65120
rect 130380 65100 130620 65120
rect 130880 65100 131120 65120
rect 131380 65100 131620 65120
rect 131880 65100 132000 65120
rect 130000 64900 132000 65100
rect 130000 64880 130120 64900
rect 130380 64880 130620 64900
rect 130880 64880 131120 64900
rect 131380 64880 131620 64900
rect 131880 64880 132000 64900
rect 130000 64620 130100 64880
rect 130400 64620 130600 64880
rect 130900 64620 131100 64880
rect 131400 64620 131600 64880
rect 131900 64620 132000 64880
rect 130000 64600 130120 64620
rect 130380 64600 130620 64620
rect 130880 64600 131120 64620
rect 131380 64600 131620 64620
rect 131880 64600 132000 64620
rect 130000 64400 132000 64600
rect 130000 64380 130120 64400
rect 130380 64380 130620 64400
rect 130880 64380 131120 64400
rect 131380 64380 131620 64400
rect 131880 64380 132000 64400
rect 130000 64120 130100 64380
rect 130400 64120 130600 64380
rect 130900 64120 131100 64380
rect 131400 64120 131600 64380
rect 131900 64120 132000 64380
rect 130000 64100 130120 64120
rect 130380 64100 130620 64120
rect 130880 64100 131120 64120
rect 131380 64100 131620 64120
rect 131880 64100 132000 64120
rect 130000 64000 132000 64100
rect 190000 65980 208000 66000
rect 190000 65910 190150 65980
rect 190350 65910 190650 65980
rect 190850 65910 191150 65980
rect 191350 65910 191650 65980
rect 191850 65910 192150 65980
rect 192350 65910 192650 65980
rect 192850 65910 193150 65980
rect 193350 65910 193650 65980
rect 193850 65910 194150 65980
rect 194350 65910 194650 65980
rect 194850 65910 195150 65980
rect 195350 65910 195650 65980
rect 195850 65910 196150 65980
rect 196350 65910 196650 65980
rect 196850 65910 197150 65980
rect 197350 65910 197650 65980
rect 197850 65910 198150 65980
rect 198350 65910 198650 65980
rect 198850 65910 199150 65980
rect 199350 65910 199650 65980
rect 199850 65910 200150 65980
rect 200350 65910 200650 65980
rect 200850 65910 201150 65980
rect 201350 65910 201650 65980
rect 201850 65910 202150 65980
rect 202350 65910 202650 65980
rect 202850 65910 203150 65980
rect 203350 65910 203650 65980
rect 203850 65910 204150 65980
rect 204350 65910 204650 65980
rect 204850 65910 205150 65980
rect 205350 65910 205650 65980
rect 205850 65910 206150 65980
rect 206350 65910 206650 65980
rect 206850 65910 207150 65980
rect 207350 65910 207650 65980
rect 207850 65910 208000 65980
rect 190000 65900 208000 65910
rect 190000 65880 190120 65900
rect 190380 65880 190620 65900
rect 190880 65880 191120 65900
rect 191380 65880 191620 65900
rect 191880 65880 192120 65900
rect 192380 65880 192620 65900
rect 192880 65880 193120 65900
rect 193380 65880 193620 65900
rect 193880 65880 194120 65900
rect 194380 65880 194620 65900
rect 194880 65880 195120 65900
rect 195380 65880 195620 65900
rect 195880 65880 196120 65900
rect 196380 65880 196620 65900
rect 196880 65880 197120 65900
rect 197380 65880 197620 65900
rect 197880 65880 198120 65900
rect 198380 65880 198620 65900
rect 198880 65880 199120 65900
rect 199380 65880 199620 65900
rect 199880 65880 200120 65900
rect 200380 65880 200620 65900
rect 200880 65880 201120 65900
rect 201380 65880 201620 65900
rect 201880 65880 202120 65900
rect 202380 65880 202620 65900
rect 202880 65880 203120 65900
rect 203380 65880 203620 65900
rect 203880 65880 204120 65900
rect 204380 65880 204620 65900
rect 204880 65880 205120 65900
rect 205380 65880 205620 65900
rect 205880 65880 206120 65900
rect 206380 65880 206620 65900
rect 206880 65880 207120 65900
rect 207380 65880 207620 65900
rect 207880 65880 208000 65900
rect 190000 65850 190100 65880
rect 190000 65650 190020 65850
rect 190090 65650 190100 65850
rect 190000 65620 190100 65650
rect 190400 65850 190600 65880
rect 190400 65650 190410 65850
rect 190480 65650 190520 65850
rect 190590 65650 190600 65850
rect 190400 65620 190600 65650
rect 190900 65850 191100 65880
rect 190900 65650 190910 65850
rect 190980 65650 191020 65850
rect 191090 65650 191100 65850
rect 190900 65620 191100 65650
rect 191400 65850 191600 65880
rect 191400 65650 191410 65850
rect 191480 65650 191520 65850
rect 191590 65650 191600 65850
rect 191400 65620 191600 65650
rect 191900 65850 192100 65880
rect 191900 65650 191910 65850
rect 191980 65650 192020 65850
rect 192090 65650 192100 65850
rect 191900 65620 192100 65650
rect 192400 65850 192600 65880
rect 192400 65650 192410 65850
rect 192480 65650 192520 65850
rect 192590 65650 192600 65850
rect 192400 65620 192600 65650
rect 192900 65850 193100 65880
rect 192900 65650 192910 65850
rect 192980 65650 193020 65850
rect 193090 65650 193100 65850
rect 192900 65620 193100 65650
rect 193400 65850 193600 65880
rect 193400 65650 193410 65850
rect 193480 65650 193520 65850
rect 193590 65650 193600 65850
rect 193400 65620 193600 65650
rect 193900 65850 194100 65880
rect 193900 65650 193910 65850
rect 193980 65650 194020 65850
rect 194090 65650 194100 65850
rect 193900 65620 194100 65650
rect 194400 65850 194600 65880
rect 194400 65650 194410 65850
rect 194480 65650 194520 65850
rect 194590 65650 194600 65850
rect 194400 65620 194600 65650
rect 194900 65850 195100 65880
rect 194900 65650 194910 65850
rect 194980 65650 195020 65850
rect 195090 65650 195100 65850
rect 194900 65620 195100 65650
rect 195400 65850 195600 65880
rect 195400 65650 195410 65850
rect 195480 65650 195520 65850
rect 195590 65650 195600 65850
rect 195400 65620 195600 65650
rect 195900 65850 196100 65880
rect 195900 65650 195910 65850
rect 195980 65650 196020 65850
rect 196090 65650 196100 65850
rect 195900 65620 196100 65650
rect 196400 65850 196600 65880
rect 196400 65650 196410 65850
rect 196480 65650 196520 65850
rect 196590 65650 196600 65850
rect 196400 65620 196600 65650
rect 196900 65850 197100 65880
rect 196900 65650 196910 65850
rect 196980 65650 197020 65850
rect 197090 65650 197100 65850
rect 196900 65620 197100 65650
rect 197400 65850 197600 65880
rect 197400 65650 197410 65850
rect 197480 65650 197520 65850
rect 197590 65650 197600 65850
rect 197400 65620 197600 65650
rect 197900 65850 198100 65880
rect 197900 65650 197910 65850
rect 197980 65650 198020 65850
rect 198090 65650 198100 65850
rect 197900 65620 198100 65650
rect 198400 65850 198600 65880
rect 198400 65650 198410 65850
rect 198480 65650 198520 65850
rect 198590 65650 198600 65850
rect 198400 65620 198600 65650
rect 198900 65850 199100 65880
rect 198900 65650 198910 65850
rect 198980 65650 199020 65850
rect 199090 65650 199100 65850
rect 198900 65620 199100 65650
rect 199400 65850 199600 65880
rect 199400 65650 199410 65850
rect 199480 65650 199520 65850
rect 199590 65650 199600 65850
rect 199400 65620 199600 65650
rect 199900 65850 200100 65880
rect 199900 65650 199910 65850
rect 199980 65650 200020 65850
rect 200090 65650 200100 65850
rect 199900 65620 200100 65650
rect 200400 65850 200600 65880
rect 200400 65650 200410 65850
rect 200480 65650 200520 65850
rect 200590 65650 200600 65850
rect 200400 65620 200600 65650
rect 200900 65850 201100 65880
rect 200900 65650 200910 65850
rect 200980 65650 201020 65850
rect 201090 65650 201100 65850
rect 200900 65620 201100 65650
rect 201400 65850 201600 65880
rect 201400 65650 201410 65850
rect 201480 65650 201520 65850
rect 201590 65650 201600 65850
rect 201400 65620 201600 65650
rect 201900 65850 202100 65880
rect 201900 65650 201910 65850
rect 201980 65650 202020 65850
rect 202090 65650 202100 65850
rect 201900 65620 202100 65650
rect 202400 65850 202600 65880
rect 202400 65650 202410 65850
rect 202480 65650 202520 65850
rect 202590 65650 202600 65850
rect 202400 65620 202600 65650
rect 202900 65850 203100 65880
rect 202900 65650 202910 65850
rect 202980 65650 203020 65850
rect 203090 65650 203100 65850
rect 202900 65620 203100 65650
rect 203400 65850 203600 65880
rect 203400 65650 203410 65850
rect 203480 65650 203520 65850
rect 203590 65650 203600 65850
rect 203400 65620 203600 65650
rect 203900 65850 204100 65880
rect 203900 65650 203910 65850
rect 203980 65650 204020 65850
rect 204090 65650 204100 65850
rect 203900 65620 204100 65650
rect 204400 65850 204600 65880
rect 204400 65650 204410 65850
rect 204480 65650 204520 65850
rect 204590 65650 204600 65850
rect 204400 65620 204600 65650
rect 204900 65850 205100 65880
rect 204900 65650 204910 65850
rect 204980 65650 205020 65850
rect 205090 65650 205100 65850
rect 204900 65620 205100 65650
rect 205400 65850 205600 65880
rect 205400 65650 205410 65850
rect 205480 65650 205520 65850
rect 205590 65650 205600 65850
rect 205400 65620 205600 65650
rect 205900 65850 206100 65880
rect 205900 65650 205910 65850
rect 205980 65650 206020 65850
rect 206090 65650 206100 65850
rect 205900 65620 206100 65650
rect 206400 65850 206600 65880
rect 206400 65650 206410 65850
rect 206480 65650 206520 65850
rect 206590 65650 206600 65850
rect 206400 65620 206600 65650
rect 206900 65850 207100 65880
rect 206900 65650 206910 65850
rect 206980 65650 207020 65850
rect 207090 65650 207100 65850
rect 206900 65620 207100 65650
rect 207400 65850 207600 65880
rect 207400 65650 207410 65850
rect 207480 65650 207520 65850
rect 207590 65650 207600 65850
rect 207400 65620 207600 65650
rect 207900 65850 208000 65880
rect 207900 65650 207910 65850
rect 207980 65650 208000 65850
rect 207900 65620 208000 65650
rect 190000 65600 190120 65620
rect 190380 65600 190620 65620
rect 190880 65600 191120 65620
rect 191380 65600 191620 65620
rect 191880 65600 192120 65620
rect 192380 65600 192620 65620
rect 192880 65600 193120 65620
rect 193380 65600 193620 65620
rect 193880 65600 194120 65620
rect 194380 65600 194620 65620
rect 194880 65600 195120 65620
rect 195380 65600 195620 65620
rect 195880 65600 196120 65620
rect 196380 65600 196620 65620
rect 196880 65600 197120 65620
rect 197380 65600 197620 65620
rect 197880 65600 198120 65620
rect 198380 65600 198620 65620
rect 198880 65600 199120 65620
rect 199380 65600 199620 65620
rect 199880 65600 200120 65620
rect 200380 65600 200620 65620
rect 200880 65600 201120 65620
rect 201380 65600 201620 65620
rect 201880 65600 202120 65620
rect 202380 65600 202620 65620
rect 202880 65600 203120 65620
rect 203380 65600 203620 65620
rect 203880 65600 204120 65620
rect 204380 65600 204620 65620
rect 204880 65600 205120 65620
rect 205380 65600 205620 65620
rect 205880 65600 206120 65620
rect 206380 65600 206620 65620
rect 206880 65600 207120 65620
rect 207380 65600 207620 65620
rect 207880 65600 208000 65620
rect 190000 65590 208000 65600
rect 190000 65520 190150 65590
rect 190350 65520 190650 65590
rect 190850 65520 191150 65590
rect 191350 65520 191650 65590
rect 191850 65520 192150 65590
rect 192350 65520 192650 65590
rect 192850 65520 193150 65590
rect 193350 65520 193650 65590
rect 193850 65520 194150 65590
rect 194350 65520 194650 65590
rect 194850 65520 195150 65590
rect 195350 65520 195650 65590
rect 195850 65520 196150 65590
rect 196350 65520 196650 65590
rect 196850 65520 197150 65590
rect 197350 65520 197650 65590
rect 197850 65520 198150 65590
rect 198350 65520 198650 65590
rect 198850 65520 199150 65590
rect 199350 65520 199650 65590
rect 199850 65520 200150 65590
rect 200350 65520 200650 65590
rect 200850 65520 201150 65590
rect 201350 65520 201650 65590
rect 201850 65520 202150 65590
rect 202350 65520 202650 65590
rect 202850 65520 203150 65590
rect 203350 65520 203650 65590
rect 203850 65520 204150 65590
rect 204350 65520 204650 65590
rect 204850 65520 205150 65590
rect 205350 65520 205650 65590
rect 205850 65520 206150 65590
rect 206350 65520 206650 65590
rect 206850 65520 207150 65590
rect 207350 65520 207650 65590
rect 207850 65520 208000 65590
rect 190000 65480 208000 65520
rect 190000 65410 190150 65480
rect 190350 65410 190650 65480
rect 190850 65410 191150 65480
rect 191350 65410 191650 65480
rect 191850 65410 192150 65480
rect 192350 65410 192650 65480
rect 192850 65410 193150 65480
rect 193350 65410 193650 65480
rect 193850 65410 194150 65480
rect 194350 65410 194650 65480
rect 194850 65410 195150 65480
rect 195350 65410 195650 65480
rect 195850 65410 196150 65480
rect 196350 65410 196650 65480
rect 196850 65410 197150 65480
rect 197350 65410 197650 65480
rect 197850 65410 198150 65480
rect 198350 65410 198650 65480
rect 198850 65410 199150 65480
rect 199350 65410 199650 65480
rect 199850 65410 200150 65480
rect 200350 65410 200650 65480
rect 200850 65410 201150 65480
rect 201350 65410 201650 65480
rect 201850 65410 202150 65480
rect 202350 65410 202650 65480
rect 202850 65410 203150 65480
rect 203350 65410 203650 65480
rect 203850 65410 204150 65480
rect 204350 65410 204650 65480
rect 204850 65410 205150 65480
rect 205350 65410 205650 65480
rect 205850 65410 206150 65480
rect 206350 65410 206650 65480
rect 206850 65410 207150 65480
rect 207350 65410 207650 65480
rect 207850 65410 208000 65480
rect 190000 65400 208000 65410
rect 190000 65380 190120 65400
rect 190380 65380 190620 65400
rect 190880 65380 191120 65400
rect 191380 65380 191620 65400
rect 191880 65380 192120 65400
rect 192380 65380 192620 65400
rect 192880 65380 193120 65400
rect 193380 65380 193620 65400
rect 193880 65380 194120 65400
rect 194380 65380 194620 65400
rect 194880 65380 195120 65400
rect 195380 65380 195620 65400
rect 195880 65380 196120 65400
rect 196380 65380 196620 65400
rect 196880 65380 197120 65400
rect 197380 65380 197620 65400
rect 197880 65380 198120 65400
rect 198380 65380 198620 65400
rect 198880 65380 199120 65400
rect 199380 65380 199620 65400
rect 199880 65380 200120 65400
rect 200380 65380 200620 65400
rect 200880 65380 201120 65400
rect 201380 65380 201620 65400
rect 201880 65380 202120 65400
rect 202380 65380 202620 65400
rect 202880 65380 203120 65400
rect 203380 65380 203620 65400
rect 203880 65380 204120 65400
rect 204380 65380 204620 65400
rect 204880 65380 205120 65400
rect 205380 65380 205620 65400
rect 205880 65380 206120 65400
rect 206380 65380 206620 65400
rect 206880 65380 207120 65400
rect 207380 65380 207620 65400
rect 207880 65380 208000 65400
rect 190000 65350 190100 65380
rect 190000 65150 190020 65350
rect 190090 65150 190100 65350
rect 190000 65120 190100 65150
rect 190400 65350 190600 65380
rect 190400 65150 190410 65350
rect 190480 65150 190520 65350
rect 190590 65150 190600 65350
rect 190400 65120 190600 65150
rect 190900 65350 191100 65380
rect 190900 65150 190910 65350
rect 190980 65150 191020 65350
rect 191090 65150 191100 65350
rect 190900 65120 191100 65150
rect 191400 65350 191600 65380
rect 191400 65150 191410 65350
rect 191480 65150 191520 65350
rect 191590 65150 191600 65350
rect 191400 65120 191600 65150
rect 191900 65350 192100 65380
rect 191900 65150 191910 65350
rect 191980 65150 192020 65350
rect 192090 65150 192100 65350
rect 191900 65120 192100 65150
rect 192400 65350 192600 65380
rect 192400 65150 192410 65350
rect 192480 65150 192520 65350
rect 192590 65150 192600 65350
rect 192400 65120 192600 65150
rect 192900 65350 193100 65380
rect 192900 65150 192910 65350
rect 192980 65150 193020 65350
rect 193090 65150 193100 65350
rect 192900 65120 193100 65150
rect 193400 65350 193600 65380
rect 193400 65150 193410 65350
rect 193480 65150 193520 65350
rect 193590 65150 193600 65350
rect 193400 65120 193600 65150
rect 193900 65350 194100 65380
rect 193900 65150 193910 65350
rect 193980 65150 194020 65350
rect 194090 65150 194100 65350
rect 193900 65120 194100 65150
rect 194400 65350 194600 65380
rect 194400 65150 194410 65350
rect 194480 65150 194520 65350
rect 194590 65150 194600 65350
rect 194400 65120 194600 65150
rect 194900 65350 195100 65380
rect 194900 65150 194910 65350
rect 194980 65150 195020 65350
rect 195090 65150 195100 65350
rect 194900 65120 195100 65150
rect 195400 65350 195600 65380
rect 195400 65150 195410 65350
rect 195480 65150 195520 65350
rect 195590 65150 195600 65350
rect 195400 65120 195600 65150
rect 195900 65350 196100 65380
rect 195900 65150 195910 65350
rect 195980 65150 196020 65350
rect 196090 65150 196100 65350
rect 195900 65120 196100 65150
rect 196400 65350 196600 65380
rect 196400 65150 196410 65350
rect 196480 65150 196520 65350
rect 196590 65150 196600 65350
rect 196400 65120 196600 65150
rect 196900 65350 197100 65380
rect 196900 65150 196910 65350
rect 196980 65150 197020 65350
rect 197090 65150 197100 65350
rect 196900 65120 197100 65150
rect 197400 65350 197600 65380
rect 197400 65150 197410 65350
rect 197480 65150 197520 65350
rect 197590 65150 197600 65350
rect 197400 65120 197600 65150
rect 197900 65350 198100 65380
rect 197900 65150 197910 65350
rect 197980 65150 198020 65350
rect 198090 65150 198100 65350
rect 197900 65120 198100 65150
rect 198400 65350 198600 65380
rect 198400 65150 198410 65350
rect 198480 65150 198520 65350
rect 198590 65150 198600 65350
rect 198400 65120 198600 65150
rect 198900 65350 199100 65380
rect 198900 65150 198910 65350
rect 198980 65150 199020 65350
rect 199090 65150 199100 65350
rect 198900 65120 199100 65150
rect 199400 65350 199600 65380
rect 199400 65150 199410 65350
rect 199480 65150 199520 65350
rect 199590 65150 199600 65350
rect 199400 65120 199600 65150
rect 199900 65350 200100 65380
rect 199900 65150 199910 65350
rect 199980 65150 200020 65350
rect 200090 65150 200100 65350
rect 199900 65120 200100 65150
rect 200400 65350 200600 65380
rect 200400 65150 200410 65350
rect 200480 65150 200520 65350
rect 200590 65150 200600 65350
rect 200400 65120 200600 65150
rect 200900 65350 201100 65380
rect 200900 65150 200910 65350
rect 200980 65150 201020 65350
rect 201090 65150 201100 65350
rect 200900 65120 201100 65150
rect 201400 65350 201600 65380
rect 201400 65150 201410 65350
rect 201480 65150 201520 65350
rect 201590 65150 201600 65350
rect 201400 65120 201600 65150
rect 201900 65350 202100 65380
rect 201900 65150 201910 65350
rect 201980 65150 202020 65350
rect 202090 65150 202100 65350
rect 201900 65120 202100 65150
rect 202400 65350 202600 65380
rect 202400 65150 202410 65350
rect 202480 65150 202520 65350
rect 202590 65150 202600 65350
rect 202400 65120 202600 65150
rect 202900 65350 203100 65380
rect 202900 65150 202910 65350
rect 202980 65150 203020 65350
rect 203090 65150 203100 65350
rect 202900 65120 203100 65150
rect 203400 65350 203600 65380
rect 203400 65150 203410 65350
rect 203480 65150 203520 65350
rect 203590 65150 203600 65350
rect 203400 65120 203600 65150
rect 203900 65350 204100 65380
rect 203900 65150 203910 65350
rect 203980 65150 204020 65350
rect 204090 65150 204100 65350
rect 203900 65120 204100 65150
rect 204400 65350 204600 65380
rect 204400 65150 204410 65350
rect 204480 65150 204520 65350
rect 204590 65150 204600 65350
rect 204400 65120 204600 65150
rect 204900 65350 205100 65380
rect 204900 65150 204910 65350
rect 204980 65150 205020 65350
rect 205090 65150 205100 65350
rect 204900 65120 205100 65150
rect 205400 65350 205600 65380
rect 205400 65150 205410 65350
rect 205480 65150 205520 65350
rect 205590 65150 205600 65350
rect 205400 65120 205600 65150
rect 205900 65350 206100 65380
rect 205900 65150 205910 65350
rect 205980 65150 206020 65350
rect 206090 65150 206100 65350
rect 205900 65120 206100 65150
rect 206400 65350 206600 65380
rect 206400 65150 206410 65350
rect 206480 65150 206520 65350
rect 206590 65150 206600 65350
rect 206400 65120 206600 65150
rect 206900 65350 207100 65380
rect 206900 65150 206910 65350
rect 206980 65150 207020 65350
rect 207090 65150 207100 65350
rect 206900 65120 207100 65150
rect 207400 65350 207600 65380
rect 207400 65150 207410 65350
rect 207480 65150 207520 65350
rect 207590 65150 207600 65350
rect 207400 65120 207600 65150
rect 207900 65350 208000 65380
rect 207900 65150 207910 65350
rect 207980 65150 208000 65350
rect 207900 65120 208000 65150
rect 190000 65100 190120 65120
rect 190380 65100 190620 65120
rect 190880 65100 191120 65120
rect 191380 65100 191620 65120
rect 191880 65100 192120 65120
rect 192380 65100 192620 65120
rect 192880 65100 193120 65120
rect 193380 65100 193620 65120
rect 193880 65100 194120 65120
rect 194380 65100 194620 65120
rect 194880 65100 195120 65120
rect 195380 65100 195620 65120
rect 195880 65100 196120 65120
rect 196380 65100 196620 65120
rect 196880 65100 197120 65120
rect 197380 65100 197620 65120
rect 197880 65100 198120 65120
rect 198380 65100 198620 65120
rect 198880 65100 199120 65120
rect 199380 65100 199620 65120
rect 199880 65100 200120 65120
rect 200380 65100 200620 65120
rect 200880 65100 201120 65120
rect 201380 65100 201620 65120
rect 201880 65100 202120 65120
rect 202380 65100 202620 65120
rect 202880 65100 203120 65120
rect 203380 65100 203620 65120
rect 203880 65100 204120 65120
rect 204380 65100 204620 65120
rect 204880 65100 205120 65120
rect 205380 65100 205620 65120
rect 205880 65100 206120 65120
rect 206380 65100 206620 65120
rect 206880 65100 207120 65120
rect 207380 65100 207620 65120
rect 207880 65100 208000 65120
rect 190000 65090 208000 65100
rect 190000 65020 190150 65090
rect 190350 65020 190650 65090
rect 190850 65020 191150 65090
rect 191350 65020 191650 65090
rect 191850 65020 192150 65090
rect 192350 65020 192650 65090
rect 192850 65020 193150 65090
rect 193350 65020 193650 65090
rect 193850 65020 194150 65090
rect 194350 65020 194650 65090
rect 194850 65020 195150 65090
rect 195350 65020 195650 65090
rect 195850 65020 196150 65090
rect 196350 65020 196650 65090
rect 196850 65020 197150 65090
rect 197350 65020 197650 65090
rect 197850 65020 198150 65090
rect 198350 65020 198650 65090
rect 198850 65020 199150 65090
rect 199350 65020 199650 65090
rect 199850 65020 200150 65090
rect 200350 65020 200650 65090
rect 200850 65020 201150 65090
rect 201350 65020 201650 65090
rect 201850 65020 202150 65090
rect 202350 65020 202650 65090
rect 202850 65020 203150 65090
rect 203350 65020 203650 65090
rect 203850 65020 204150 65090
rect 204350 65020 204650 65090
rect 204850 65020 205150 65090
rect 205350 65020 205650 65090
rect 205850 65020 206150 65090
rect 206350 65020 206650 65090
rect 206850 65020 207150 65090
rect 207350 65020 207650 65090
rect 207850 65020 208000 65090
rect 190000 64980 208000 65020
rect 190000 64910 190150 64980
rect 190350 64910 190650 64980
rect 190850 64910 191150 64980
rect 191350 64910 191650 64980
rect 191850 64910 192150 64980
rect 192350 64910 192650 64980
rect 192850 64910 193150 64980
rect 193350 64910 193650 64980
rect 193850 64910 194150 64980
rect 194350 64910 194650 64980
rect 194850 64910 195150 64980
rect 195350 64910 195650 64980
rect 195850 64910 196150 64980
rect 196350 64910 196650 64980
rect 196850 64910 197150 64980
rect 197350 64910 197650 64980
rect 197850 64910 198150 64980
rect 198350 64910 198650 64980
rect 198850 64910 199150 64980
rect 199350 64910 199650 64980
rect 199850 64910 200150 64980
rect 200350 64910 200650 64980
rect 200850 64910 201150 64980
rect 201350 64910 201650 64980
rect 201850 64910 202150 64980
rect 202350 64910 202650 64980
rect 202850 64910 203150 64980
rect 203350 64910 203650 64980
rect 203850 64910 204150 64980
rect 204350 64910 204650 64980
rect 204850 64910 205150 64980
rect 205350 64910 205650 64980
rect 205850 64910 206150 64980
rect 206350 64910 206650 64980
rect 206850 64910 207150 64980
rect 207350 64910 207650 64980
rect 207850 64910 208000 64980
rect 190000 64900 208000 64910
rect 190000 64880 190120 64900
rect 190380 64880 190620 64900
rect 190880 64880 191120 64900
rect 191380 64880 191620 64900
rect 191880 64880 192120 64900
rect 192380 64880 192620 64900
rect 192880 64880 193120 64900
rect 193380 64880 193620 64900
rect 193880 64880 194120 64900
rect 194380 64880 194620 64900
rect 194880 64880 195120 64900
rect 195380 64880 195620 64900
rect 195880 64880 196120 64900
rect 196380 64880 196620 64900
rect 196880 64880 197120 64900
rect 197380 64880 197620 64900
rect 197880 64880 198120 64900
rect 198380 64880 198620 64900
rect 198880 64880 199120 64900
rect 199380 64880 199620 64900
rect 199880 64880 200120 64900
rect 200380 64880 200620 64900
rect 200880 64880 201120 64900
rect 201380 64880 201620 64900
rect 201880 64880 202120 64900
rect 202380 64880 202620 64900
rect 202880 64880 203120 64900
rect 203380 64880 203620 64900
rect 203880 64880 204120 64900
rect 204380 64880 204620 64900
rect 204880 64880 205120 64900
rect 205380 64880 205620 64900
rect 205880 64880 206120 64900
rect 206380 64880 206620 64900
rect 206880 64880 207120 64900
rect 207380 64880 207620 64900
rect 207880 64880 208000 64900
rect 190000 64850 190100 64880
rect 190000 64650 190020 64850
rect 190090 64650 190100 64850
rect 190000 64620 190100 64650
rect 190400 64850 190600 64880
rect 190400 64650 190410 64850
rect 190480 64650 190520 64850
rect 190590 64650 190600 64850
rect 190400 64620 190600 64650
rect 190900 64850 191100 64880
rect 190900 64650 190910 64850
rect 190980 64650 191020 64850
rect 191090 64650 191100 64850
rect 190900 64620 191100 64650
rect 191400 64850 191600 64880
rect 191400 64650 191410 64850
rect 191480 64650 191520 64850
rect 191590 64650 191600 64850
rect 191400 64620 191600 64650
rect 191900 64850 192100 64880
rect 191900 64650 191910 64850
rect 191980 64650 192020 64850
rect 192090 64650 192100 64850
rect 191900 64620 192100 64650
rect 192400 64850 192600 64880
rect 192400 64650 192410 64850
rect 192480 64650 192520 64850
rect 192590 64650 192600 64850
rect 192400 64620 192600 64650
rect 192900 64850 193100 64880
rect 192900 64650 192910 64850
rect 192980 64650 193020 64850
rect 193090 64650 193100 64850
rect 192900 64620 193100 64650
rect 193400 64850 193600 64880
rect 193400 64650 193410 64850
rect 193480 64650 193520 64850
rect 193590 64650 193600 64850
rect 193400 64620 193600 64650
rect 193900 64850 194100 64880
rect 193900 64650 193910 64850
rect 193980 64650 194020 64850
rect 194090 64650 194100 64850
rect 193900 64620 194100 64650
rect 194400 64850 194600 64880
rect 194400 64650 194410 64850
rect 194480 64650 194520 64850
rect 194590 64650 194600 64850
rect 194400 64620 194600 64650
rect 194900 64850 195100 64880
rect 194900 64650 194910 64850
rect 194980 64650 195020 64850
rect 195090 64650 195100 64850
rect 194900 64620 195100 64650
rect 195400 64850 195600 64880
rect 195400 64650 195410 64850
rect 195480 64650 195520 64850
rect 195590 64650 195600 64850
rect 195400 64620 195600 64650
rect 195900 64850 196100 64880
rect 195900 64650 195910 64850
rect 195980 64650 196020 64850
rect 196090 64650 196100 64850
rect 195900 64620 196100 64650
rect 196400 64850 196600 64880
rect 196400 64650 196410 64850
rect 196480 64650 196520 64850
rect 196590 64650 196600 64850
rect 196400 64620 196600 64650
rect 196900 64850 197100 64880
rect 196900 64650 196910 64850
rect 196980 64650 197020 64850
rect 197090 64650 197100 64850
rect 196900 64620 197100 64650
rect 197400 64850 197600 64880
rect 197400 64650 197410 64850
rect 197480 64650 197520 64850
rect 197590 64650 197600 64850
rect 197400 64620 197600 64650
rect 197900 64850 198100 64880
rect 197900 64650 197910 64850
rect 197980 64650 198020 64850
rect 198090 64650 198100 64850
rect 197900 64620 198100 64650
rect 198400 64850 198600 64880
rect 198400 64650 198410 64850
rect 198480 64650 198520 64850
rect 198590 64650 198600 64850
rect 198400 64620 198600 64650
rect 198900 64850 199100 64880
rect 198900 64650 198910 64850
rect 198980 64650 199020 64850
rect 199090 64650 199100 64850
rect 198900 64620 199100 64650
rect 199400 64850 199600 64880
rect 199400 64650 199410 64850
rect 199480 64650 199520 64850
rect 199590 64650 199600 64850
rect 199400 64620 199600 64650
rect 199900 64850 200100 64880
rect 199900 64650 199910 64850
rect 199980 64650 200020 64850
rect 200090 64650 200100 64850
rect 199900 64620 200100 64650
rect 200400 64850 200600 64880
rect 200400 64650 200410 64850
rect 200480 64650 200520 64850
rect 200590 64650 200600 64850
rect 200400 64620 200600 64650
rect 200900 64850 201100 64880
rect 200900 64650 200910 64850
rect 200980 64650 201020 64850
rect 201090 64650 201100 64850
rect 200900 64620 201100 64650
rect 201400 64850 201600 64880
rect 201400 64650 201410 64850
rect 201480 64650 201520 64850
rect 201590 64650 201600 64850
rect 201400 64620 201600 64650
rect 201900 64850 202100 64880
rect 201900 64650 201910 64850
rect 201980 64650 202020 64850
rect 202090 64650 202100 64850
rect 201900 64620 202100 64650
rect 202400 64850 202600 64880
rect 202400 64650 202410 64850
rect 202480 64650 202520 64850
rect 202590 64650 202600 64850
rect 202400 64620 202600 64650
rect 202900 64850 203100 64880
rect 202900 64650 202910 64850
rect 202980 64650 203020 64850
rect 203090 64650 203100 64850
rect 202900 64620 203100 64650
rect 203400 64850 203600 64880
rect 203400 64650 203410 64850
rect 203480 64650 203520 64850
rect 203590 64650 203600 64850
rect 203400 64620 203600 64650
rect 203900 64850 204100 64880
rect 203900 64650 203910 64850
rect 203980 64650 204020 64850
rect 204090 64650 204100 64850
rect 203900 64620 204100 64650
rect 204400 64850 204600 64880
rect 204400 64650 204410 64850
rect 204480 64650 204520 64850
rect 204590 64650 204600 64850
rect 204400 64620 204600 64650
rect 204900 64850 205100 64880
rect 204900 64650 204910 64850
rect 204980 64650 205020 64850
rect 205090 64650 205100 64850
rect 204900 64620 205100 64650
rect 205400 64850 205600 64880
rect 205400 64650 205410 64850
rect 205480 64650 205520 64850
rect 205590 64650 205600 64850
rect 205400 64620 205600 64650
rect 205900 64850 206100 64880
rect 205900 64650 205910 64850
rect 205980 64650 206020 64850
rect 206090 64650 206100 64850
rect 205900 64620 206100 64650
rect 206400 64850 206600 64880
rect 206400 64650 206410 64850
rect 206480 64650 206520 64850
rect 206590 64650 206600 64850
rect 206400 64620 206600 64650
rect 206900 64850 207100 64880
rect 206900 64650 206910 64850
rect 206980 64650 207020 64850
rect 207090 64650 207100 64850
rect 206900 64620 207100 64650
rect 207400 64850 207600 64880
rect 207400 64650 207410 64850
rect 207480 64650 207520 64850
rect 207590 64650 207600 64850
rect 207400 64620 207600 64650
rect 207900 64850 208000 64880
rect 207900 64650 207910 64850
rect 207980 64650 208000 64850
rect 207900 64620 208000 64650
rect 190000 64600 190120 64620
rect 190380 64600 190620 64620
rect 190880 64600 191120 64620
rect 191380 64600 191620 64620
rect 191880 64600 192120 64620
rect 192380 64600 192620 64620
rect 192880 64600 193120 64620
rect 193380 64600 193620 64620
rect 193880 64600 194120 64620
rect 194380 64600 194620 64620
rect 194880 64600 195120 64620
rect 195380 64600 195620 64620
rect 195880 64600 196120 64620
rect 196380 64600 196620 64620
rect 196880 64600 197120 64620
rect 197380 64600 197620 64620
rect 197880 64600 198120 64620
rect 198380 64600 198620 64620
rect 198880 64600 199120 64620
rect 199380 64600 199620 64620
rect 199880 64600 200120 64620
rect 200380 64600 200620 64620
rect 200880 64600 201120 64620
rect 201380 64600 201620 64620
rect 201880 64600 202120 64620
rect 202380 64600 202620 64620
rect 202880 64600 203120 64620
rect 203380 64600 203620 64620
rect 203880 64600 204120 64620
rect 204380 64600 204620 64620
rect 204880 64600 205120 64620
rect 205380 64600 205620 64620
rect 205880 64600 206120 64620
rect 206380 64600 206620 64620
rect 206880 64600 207120 64620
rect 207380 64600 207620 64620
rect 207880 64600 208000 64620
rect 190000 64590 208000 64600
rect 190000 64520 190150 64590
rect 190350 64520 190650 64590
rect 190850 64520 191150 64590
rect 191350 64520 191650 64590
rect 191850 64520 192150 64590
rect 192350 64520 192650 64590
rect 192850 64520 193150 64590
rect 193350 64520 193650 64590
rect 193850 64520 194150 64590
rect 194350 64520 194650 64590
rect 194850 64520 195150 64590
rect 195350 64520 195650 64590
rect 195850 64520 196150 64590
rect 196350 64520 196650 64590
rect 196850 64520 197150 64590
rect 197350 64520 197650 64590
rect 197850 64520 198150 64590
rect 198350 64520 198650 64590
rect 198850 64520 199150 64590
rect 199350 64520 199650 64590
rect 199850 64520 200150 64590
rect 200350 64520 200650 64590
rect 200850 64520 201150 64590
rect 201350 64520 201650 64590
rect 201850 64520 202150 64590
rect 202350 64520 202650 64590
rect 202850 64520 203150 64590
rect 203350 64520 203650 64590
rect 203850 64520 204150 64590
rect 204350 64520 204650 64590
rect 204850 64520 205150 64590
rect 205350 64520 205650 64590
rect 205850 64520 206150 64590
rect 206350 64520 206650 64590
rect 206850 64520 207150 64590
rect 207350 64520 207650 64590
rect 207850 64520 208000 64590
rect 190000 64480 208000 64520
rect 190000 64410 190150 64480
rect 190350 64410 190650 64480
rect 190850 64410 191150 64480
rect 191350 64410 191650 64480
rect 191850 64410 192150 64480
rect 192350 64410 192650 64480
rect 192850 64410 193150 64480
rect 193350 64410 193650 64480
rect 193850 64410 194150 64480
rect 194350 64410 194650 64480
rect 194850 64410 195150 64480
rect 195350 64410 195650 64480
rect 195850 64410 196150 64480
rect 196350 64410 196650 64480
rect 196850 64410 197150 64480
rect 197350 64410 197650 64480
rect 197850 64410 198150 64480
rect 198350 64410 198650 64480
rect 198850 64410 199150 64480
rect 199350 64410 199650 64480
rect 199850 64410 200150 64480
rect 200350 64410 200650 64480
rect 200850 64410 201150 64480
rect 201350 64410 201650 64480
rect 201850 64410 202150 64480
rect 202350 64410 202650 64480
rect 202850 64410 203150 64480
rect 203350 64410 203650 64480
rect 203850 64410 204150 64480
rect 204350 64410 204650 64480
rect 204850 64410 205150 64480
rect 205350 64410 205650 64480
rect 205850 64410 206150 64480
rect 206350 64410 206650 64480
rect 206850 64410 207150 64480
rect 207350 64410 207650 64480
rect 207850 64410 208000 64480
rect 190000 64400 208000 64410
rect 190000 64380 190120 64400
rect 190380 64380 190620 64400
rect 190880 64380 191120 64400
rect 191380 64380 191620 64400
rect 191880 64380 192120 64400
rect 192380 64380 192620 64400
rect 192880 64380 193120 64400
rect 193380 64380 193620 64400
rect 193880 64380 194120 64400
rect 194380 64380 194620 64400
rect 194880 64380 195120 64400
rect 195380 64380 195620 64400
rect 195880 64380 196120 64400
rect 196380 64380 196620 64400
rect 196880 64380 197120 64400
rect 197380 64380 197620 64400
rect 197880 64380 198120 64400
rect 198380 64380 198620 64400
rect 198880 64380 199120 64400
rect 199380 64380 199620 64400
rect 199880 64380 200120 64400
rect 200380 64380 200620 64400
rect 200880 64380 201120 64400
rect 201380 64380 201620 64400
rect 201880 64380 202120 64400
rect 202380 64380 202620 64400
rect 202880 64380 203120 64400
rect 203380 64380 203620 64400
rect 203880 64380 204120 64400
rect 204380 64380 204620 64400
rect 204880 64380 205120 64400
rect 205380 64380 205620 64400
rect 205880 64380 206120 64400
rect 206380 64380 206620 64400
rect 206880 64380 207120 64400
rect 207380 64380 207620 64400
rect 207880 64380 208000 64400
rect 190000 64350 190100 64380
rect 190000 64150 190020 64350
rect 190090 64150 190100 64350
rect 190000 64120 190100 64150
rect 190400 64350 190600 64380
rect 190400 64150 190410 64350
rect 190480 64150 190520 64350
rect 190590 64150 190600 64350
rect 190400 64120 190600 64150
rect 190900 64350 191100 64380
rect 190900 64150 190910 64350
rect 190980 64150 191020 64350
rect 191090 64150 191100 64350
rect 190900 64120 191100 64150
rect 191400 64350 191600 64380
rect 191400 64150 191410 64350
rect 191480 64150 191520 64350
rect 191590 64150 191600 64350
rect 191400 64120 191600 64150
rect 191900 64350 192100 64380
rect 191900 64150 191910 64350
rect 191980 64150 192020 64350
rect 192090 64150 192100 64350
rect 191900 64120 192100 64150
rect 192400 64350 192600 64380
rect 192400 64150 192410 64350
rect 192480 64150 192520 64350
rect 192590 64150 192600 64350
rect 192400 64120 192600 64150
rect 192900 64350 193100 64380
rect 192900 64150 192910 64350
rect 192980 64150 193020 64350
rect 193090 64150 193100 64350
rect 192900 64120 193100 64150
rect 193400 64350 193600 64380
rect 193400 64150 193410 64350
rect 193480 64150 193520 64350
rect 193590 64150 193600 64350
rect 193400 64120 193600 64150
rect 193900 64350 194100 64380
rect 193900 64150 193910 64350
rect 193980 64150 194020 64350
rect 194090 64150 194100 64350
rect 193900 64120 194100 64150
rect 194400 64350 194600 64380
rect 194400 64150 194410 64350
rect 194480 64150 194520 64350
rect 194590 64150 194600 64350
rect 194400 64120 194600 64150
rect 194900 64350 195100 64380
rect 194900 64150 194910 64350
rect 194980 64150 195020 64350
rect 195090 64150 195100 64350
rect 194900 64120 195100 64150
rect 195400 64350 195600 64380
rect 195400 64150 195410 64350
rect 195480 64150 195520 64350
rect 195590 64150 195600 64350
rect 195400 64120 195600 64150
rect 195900 64350 196100 64380
rect 195900 64150 195910 64350
rect 195980 64150 196020 64350
rect 196090 64150 196100 64350
rect 195900 64120 196100 64150
rect 196400 64350 196600 64380
rect 196400 64150 196410 64350
rect 196480 64150 196520 64350
rect 196590 64150 196600 64350
rect 196400 64120 196600 64150
rect 196900 64350 197100 64380
rect 196900 64150 196910 64350
rect 196980 64150 197020 64350
rect 197090 64150 197100 64350
rect 196900 64120 197100 64150
rect 197400 64350 197600 64380
rect 197400 64150 197410 64350
rect 197480 64150 197520 64350
rect 197590 64150 197600 64350
rect 197400 64120 197600 64150
rect 197900 64350 198100 64380
rect 197900 64150 197910 64350
rect 197980 64150 198020 64350
rect 198090 64150 198100 64350
rect 197900 64120 198100 64150
rect 198400 64350 198600 64380
rect 198400 64150 198410 64350
rect 198480 64150 198520 64350
rect 198590 64150 198600 64350
rect 198400 64120 198600 64150
rect 198900 64350 199100 64380
rect 198900 64150 198910 64350
rect 198980 64150 199020 64350
rect 199090 64150 199100 64350
rect 198900 64120 199100 64150
rect 199400 64350 199600 64380
rect 199400 64150 199410 64350
rect 199480 64150 199520 64350
rect 199590 64150 199600 64350
rect 199400 64120 199600 64150
rect 199900 64350 200100 64380
rect 199900 64150 199910 64350
rect 199980 64150 200020 64350
rect 200090 64150 200100 64350
rect 199900 64120 200100 64150
rect 200400 64350 200600 64380
rect 200400 64150 200410 64350
rect 200480 64150 200520 64350
rect 200590 64150 200600 64350
rect 200400 64120 200600 64150
rect 200900 64350 201100 64380
rect 200900 64150 200910 64350
rect 200980 64150 201020 64350
rect 201090 64150 201100 64350
rect 200900 64120 201100 64150
rect 201400 64350 201600 64380
rect 201400 64150 201410 64350
rect 201480 64150 201520 64350
rect 201590 64150 201600 64350
rect 201400 64120 201600 64150
rect 201900 64350 202100 64380
rect 201900 64150 201910 64350
rect 201980 64150 202020 64350
rect 202090 64150 202100 64350
rect 201900 64120 202100 64150
rect 202400 64350 202600 64380
rect 202400 64150 202410 64350
rect 202480 64150 202520 64350
rect 202590 64150 202600 64350
rect 202400 64120 202600 64150
rect 202900 64350 203100 64380
rect 202900 64150 202910 64350
rect 202980 64150 203020 64350
rect 203090 64150 203100 64350
rect 202900 64120 203100 64150
rect 203400 64350 203600 64380
rect 203400 64150 203410 64350
rect 203480 64150 203520 64350
rect 203590 64150 203600 64350
rect 203400 64120 203600 64150
rect 203900 64350 204100 64380
rect 203900 64150 203910 64350
rect 203980 64150 204020 64350
rect 204090 64150 204100 64350
rect 203900 64120 204100 64150
rect 204400 64350 204600 64380
rect 204400 64150 204410 64350
rect 204480 64150 204520 64350
rect 204590 64150 204600 64350
rect 204400 64120 204600 64150
rect 204900 64350 205100 64380
rect 204900 64150 204910 64350
rect 204980 64150 205020 64350
rect 205090 64150 205100 64350
rect 204900 64120 205100 64150
rect 205400 64350 205600 64380
rect 205400 64150 205410 64350
rect 205480 64150 205520 64350
rect 205590 64150 205600 64350
rect 205400 64120 205600 64150
rect 205900 64350 206100 64380
rect 205900 64150 205910 64350
rect 205980 64150 206020 64350
rect 206090 64150 206100 64350
rect 205900 64120 206100 64150
rect 206400 64350 206600 64380
rect 206400 64150 206410 64350
rect 206480 64150 206520 64350
rect 206590 64150 206600 64350
rect 206400 64120 206600 64150
rect 206900 64350 207100 64380
rect 206900 64150 206910 64350
rect 206980 64150 207020 64350
rect 207090 64150 207100 64350
rect 206900 64120 207100 64150
rect 207400 64350 207600 64380
rect 207400 64150 207410 64350
rect 207480 64150 207520 64350
rect 207590 64150 207600 64350
rect 207400 64120 207600 64150
rect 207900 64350 208000 64380
rect 207900 64150 207910 64350
rect 207980 64150 208000 64350
rect 207900 64120 208000 64150
rect 190000 64100 190120 64120
rect 190380 64100 190620 64120
rect 190880 64100 191120 64120
rect 191380 64100 191620 64120
rect 191880 64100 192120 64120
rect 192380 64100 192620 64120
rect 192880 64100 193120 64120
rect 193380 64100 193620 64120
rect 193880 64100 194120 64120
rect 194380 64100 194620 64120
rect 194880 64100 195120 64120
rect 195380 64100 195620 64120
rect 195880 64100 196120 64120
rect 196380 64100 196620 64120
rect 196880 64100 197120 64120
rect 197380 64100 197620 64120
rect 197880 64100 198120 64120
rect 198380 64100 198620 64120
rect 198880 64100 199120 64120
rect 199380 64100 199620 64120
rect 199880 64100 200120 64120
rect 200380 64100 200620 64120
rect 200880 64100 201120 64120
rect 201380 64100 201620 64120
rect 201880 64100 202120 64120
rect 202380 64100 202620 64120
rect 202880 64100 203120 64120
rect 203380 64100 203620 64120
rect 203880 64100 204120 64120
rect 204380 64100 204620 64120
rect 204880 64100 205120 64120
rect 205380 64100 205620 64120
rect 205880 64100 206120 64120
rect 206380 64100 206620 64120
rect 206880 64100 207120 64120
rect 207380 64100 207620 64120
rect 207880 64100 208000 64120
rect 190000 64090 208000 64100
rect 190000 64020 190150 64090
rect 190350 64020 190650 64090
rect 190850 64020 191150 64090
rect 191350 64020 191650 64090
rect 191850 64020 192150 64090
rect 192350 64020 192650 64090
rect 192850 64020 193150 64090
rect 193350 64020 193650 64090
rect 193850 64020 194150 64090
rect 194350 64020 194650 64090
rect 194850 64020 195150 64090
rect 195350 64020 195650 64090
rect 195850 64020 196150 64090
rect 196350 64020 196650 64090
rect 196850 64020 197150 64090
rect 197350 64020 197650 64090
rect 197850 64020 198150 64090
rect 198350 64020 198650 64090
rect 198850 64020 199150 64090
rect 199350 64020 199650 64090
rect 199850 64020 200150 64090
rect 200350 64020 200650 64090
rect 200850 64020 201150 64090
rect 201350 64020 201650 64090
rect 201850 64020 202150 64090
rect 202350 64020 202650 64090
rect 202850 64020 203150 64090
rect 203350 64020 203650 64090
rect 203850 64020 204150 64090
rect 204350 64020 204650 64090
rect 204850 64020 205150 64090
rect 205350 64020 205650 64090
rect 205850 64020 206150 64090
rect 206350 64020 206650 64090
rect 206850 64020 207150 64090
rect 207350 64020 207650 64090
rect 207850 64020 208000 64090
rect 190000 64000 208000 64020
rect 132000 63900 135000 64000
rect 132000 63880 132120 63900
rect 132380 63880 132620 63900
rect 132880 63880 133120 63900
rect 133380 63880 133620 63900
rect 133880 63880 134120 63900
rect 134380 63880 134620 63900
rect 134880 63880 135000 63900
rect 132000 63620 132100 63880
rect 132400 63620 132600 63880
rect 132900 63620 133100 63880
rect 133400 63620 133600 63880
rect 133900 63620 134100 63880
rect 134400 63620 134600 63880
rect 134900 63620 135000 63880
rect 132000 63600 132120 63620
rect 132380 63600 132620 63620
rect 132880 63600 133120 63620
rect 133380 63600 133620 63620
rect 133880 63600 134120 63620
rect 134380 63600 134620 63620
rect 134880 63600 135000 63620
rect 132000 63400 135000 63600
rect 132000 63380 132120 63400
rect 132380 63380 132620 63400
rect 132880 63380 133120 63400
rect 133380 63380 133620 63400
rect 133880 63380 134120 63400
rect 134380 63380 134620 63400
rect 134880 63380 135000 63400
rect 132000 63120 132100 63380
rect 132400 63120 132600 63380
rect 132900 63120 133100 63380
rect 133400 63120 133600 63380
rect 133900 63120 134100 63380
rect 134400 63120 134600 63380
rect 134900 63120 135000 63380
rect 132000 63100 132120 63120
rect 132380 63100 132620 63120
rect 132880 63100 133120 63120
rect 133380 63100 133620 63120
rect 133880 63100 134120 63120
rect 134380 63100 134620 63120
rect 134880 63100 135000 63120
rect 132000 62900 135000 63100
rect 132000 62880 132120 62900
rect 132380 62880 132620 62900
rect 132880 62880 133120 62900
rect 133380 62880 133620 62900
rect 133880 62880 134120 62900
rect 134380 62880 134620 62900
rect 134880 62880 135000 62900
rect 132000 62620 132100 62880
rect 132400 62620 132600 62880
rect 132900 62620 133100 62880
rect 133400 62620 133600 62880
rect 133900 62620 134100 62880
rect 134400 62620 134600 62880
rect 134900 62620 135000 62880
rect 132000 62600 132120 62620
rect 132380 62600 132620 62620
rect 132880 62600 133120 62620
rect 133380 62600 133620 62620
rect 133880 62600 134120 62620
rect 134380 62600 134620 62620
rect 134880 62600 135000 62620
rect 132000 62400 135000 62600
rect 132000 62380 132120 62400
rect 132380 62380 132620 62400
rect 132880 62380 133120 62400
rect 133380 62380 133620 62400
rect 133880 62380 134120 62400
rect 134380 62380 134620 62400
rect 134880 62380 135000 62400
rect 132000 62120 132100 62380
rect 132400 62120 132600 62380
rect 132900 62120 133100 62380
rect 133400 62120 133600 62380
rect 133900 62120 134100 62380
rect 134400 62120 134600 62380
rect 134900 62120 135000 62380
rect 132000 62100 132120 62120
rect 132380 62100 132620 62120
rect 132880 62100 133120 62120
rect 133380 62100 133620 62120
rect 133880 62100 134120 62120
rect 134380 62100 134620 62120
rect 134880 62100 135000 62120
rect 132000 61900 135000 62100
rect 132000 61880 132120 61900
rect 132380 61880 132620 61900
rect 132880 61880 133120 61900
rect 133380 61880 133620 61900
rect 133880 61880 134120 61900
rect 134380 61880 134620 61900
rect 134880 61880 135000 61900
rect 132000 61620 132100 61880
rect 132400 61620 132600 61880
rect 132900 61620 133100 61880
rect 133400 61620 133600 61880
rect 133900 61620 134100 61880
rect 134400 61620 134600 61880
rect 134900 61620 135000 61880
rect 132000 61600 132120 61620
rect 132380 61600 132620 61620
rect 132880 61600 133120 61620
rect 133380 61600 133620 61620
rect 133880 61600 134120 61620
rect 134380 61600 134620 61620
rect 134880 61600 135000 61620
rect 132000 61400 135000 61600
rect 132000 61380 132120 61400
rect 132380 61380 132620 61400
rect 132880 61380 133120 61400
rect 133380 61380 133620 61400
rect 133880 61380 134120 61400
rect 134380 61380 134620 61400
rect 134880 61380 135000 61400
rect 132000 61120 132100 61380
rect 132400 61120 132600 61380
rect 132900 61120 133100 61380
rect 133400 61120 133600 61380
rect 133900 61120 134100 61380
rect 134400 61120 134600 61380
rect 134900 61120 135000 61380
rect 132000 61100 132120 61120
rect 132380 61100 132620 61120
rect 132880 61100 133120 61120
rect 133380 61100 133620 61120
rect 133880 61100 134120 61120
rect 134380 61100 134620 61120
rect 134880 61100 135000 61120
rect 132000 60900 135000 61100
rect 132000 60880 132120 60900
rect 132380 60880 132620 60900
rect 132880 60880 133120 60900
rect 133380 60880 133620 60900
rect 133880 60880 134120 60900
rect 134380 60880 134620 60900
rect 134880 60880 135000 60900
rect 132000 60620 132100 60880
rect 132400 60620 132600 60880
rect 132900 60620 133100 60880
rect 133400 60620 133600 60880
rect 133900 60620 134100 60880
rect 134400 60620 134600 60880
rect 134900 60620 135000 60880
rect 132000 60600 132120 60620
rect 132380 60600 132620 60620
rect 132880 60600 133120 60620
rect 133380 60600 133620 60620
rect 133880 60600 134120 60620
rect 134380 60600 134620 60620
rect 134880 60600 135000 60620
rect 132000 60400 135000 60600
rect 132000 60380 132120 60400
rect 132380 60380 132620 60400
rect 132880 60380 133120 60400
rect 133380 60380 133620 60400
rect 133880 60380 134120 60400
rect 134380 60380 134620 60400
rect 134880 60380 135000 60400
rect 132000 60120 132100 60380
rect 132400 60120 132600 60380
rect 132900 60120 133100 60380
rect 133400 60120 133600 60380
rect 133900 60120 134100 60380
rect 134400 60120 134600 60380
rect 134900 60120 135000 60380
rect 132000 60100 132120 60120
rect 132380 60100 132620 60120
rect 132880 60100 133120 60120
rect 133380 60100 133620 60120
rect 133880 60100 134120 60120
rect 134380 60100 134620 60120
rect 134880 60100 135000 60120
rect 132000 59900 135000 60100
rect 132000 59880 132120 59900
rect 132380 59880 132620 59900
rect 132880 59880 133120 59900
rect 133380 59880 133620 59900
rect 133880 59880 134120 59900
rect 134380 59880 134620 59900
rect 134880 59880 135000 59900
rect 132000 59620 132100 59880
rect 132400 59620 132600 59880
rect 132900 59620 133100 59880
rect 133400 59620 133600 59880
rect 133900 59620 134100 59880
rect 134400 59620 134600 59880
rect 134900 59620 135000 59880
rect 132000 59600 132120 59620
rect 132380 59600 132620 59620
rect 132880 59600 133120 59620
rect 133380 59600 133620 59620
rect 133880 59600 134120 59620
rect 134380 59600 134620 59620
rect 134880 59600 135000 59620
rect 132000 59400 135000 59600
rect 132000 59380 132120 59400
rect 132380 59380 132620 59400
rect 132880 59380 133120 59400
rect 133380 59380 133620 59400
rect 133880 59380 134120 59400
rect 134380 59380 134620 59400
rect 134880 59380 135000 59400
rect 132000 59120 132100 59380
rect 132400 59120 132600 59380
rect 132900 59120 133100 59380
rect 133400 59120 133600 59380
rect 133900 59120 134100 59380
rect 134400 59120 134600 59380
rect 134900 59120 135000 59380
rect 132000 59100 132120 59120
rect 132380 59100 132620 59120
rect 132880 59100 133120 59120
rect 133380 59100 133620 59120
rect 133880 59100 134120 59120
rect 134380 59100 134620 59120
rect 134880 59100 135000 59120
rect 132000 58900 135000 59100
rect 132000 58880 132120 58900
rect 132380 58880 132620 58900
rect 132880 58880 133120 58900
rect 133380 58880 133620 58900
rect 133880 58880 134120 58900
rect 134380 58880 134620 58900
rect 134880 58880 135000 58900
rect 132000 58620 132100 58880
rect 132400 58620 132600 58880
rect 132900 58620 133100 58880
rect 133400 58620 133600 58880
rect 133900 58620 134100 58880
rect 134400 58620 134600 58880
rect 134900 58620 135000 58880
rect 132000 58600 132120 58620
rect 132380 58600 132620 58620
rect 132880 58600 133120 58620
rect 133380 58600 133620 58620
rect 133880 58600 134120 58620
rect 134380 58600 134620 58620
rect 134880 58600 135000 58620
rect 132000 58400 135000 58600
rect 132000 58380 132120 58400
rect 132380 58380 132620 58400
rect 132880 58380 133120 58400
rect 133380 58380 133620 58400
rect 133880 58380 134120 58400
rect 134380 58380 134620 58400
rect 134880 58380 135000 58400
rect 132000 58120 132100 58380
rect 132400 58120 132600 58380
rect 132900 58120 133100 58380
rect 133400 58120 133600 58380
rect 133900 58120 134100 58380
rect 134400 58120 134600 58380
rect 134900 58120 135000 58380
rect 132000 58100 132120 58120
rect 132380 58100 132620 58120
rect 132880 58100 133120 58120
rect 133380 58100 133620 58120
rect 133880 58100 134120 58120
rect 134380 58100 134620 58120
rect 134880 58100 135000 58120
rect 132000 57900 135000 58100
rect 132000 57880 132120 57900
rect 132380 57880 132620 57900
rect 132880 57880 133120 57900
rect 133380 57880 133620 57900
rect 133880 57880 134120 57900
rect 134380 57880 134620 57900
rect 134880 57880 135000 57900
rect 132000 57620 132100 57880
rect 132400 57620 132600 57880
rect 132900 57620 133100 57880
rect 133400 57620 133600 57880
rect 133900 57620 134100 57880
rect 134400 57620 134600 57880
rect 134900 57620 135000 57880
rect 132000 57600 132120 57620
rect 132380 57600 132620 57620
rect 132880 57600 133120 57620
rect 133380 57600 133620 57620
rect 133880 57600 134120 57620
rect 134380 57600 134620 57620
rect 134880 57600 135000 57620
rect 132000 57400 135000 57600
rect 132000 57380 132120 57400
rect 132380 57380 132620 57400
rect 132880 57380 133120 57400
rect 133380 57380 133620 57400
rect 133880 57380 134120 57400
rect 134380 57380 134620 57400
rect 134880 57380 135000 57400
rect 132000 57120 132100 57380
rect 132400 57120 132600 57380
rect 132900 57120 133100 57380
rect 133400 57120 133600 57380
rect 133900 57120 134100 57380
rect 134400 57120 134600 57380
rect 134900 57120 135000 57380
rect 132000 57100 132120 57120
rect 132380 57100 132620 57120
rect 132880 57100 133120 57120
rect 133380 57100 133620 57120
rect 133880 57100 134120 57120
rect 134380 57100 134620 57120
rect 134880 57100 135000 57120
rect 132000 56900 135000 57100
rect 132000 56880 132120 56900
rect 132380 56880 132620 56900
rect 132880 56880 133120 56900
rect 133380 56880 133620 56900
rect 133880 56880 134120 56900
rect 134380 56880 134620 56900
rect 134880 56880 135000 56900
rect 132000 56620 132100 56880
rect 132400 56620 132600 56880
rect 132900 56620 133100 56880
rect 133400 56620 133600 56880
rect 133900 56620 134100 56880
rect 134400 56620 134600 56880
rect 134900 56620 135000 56880
rect 132000 56600 132120 56620
rect 132380 56600 132620 56620
rect 132880 56600 133120 56620
rect 133380 56600 133620 56620
rect 133880 56600 134120 56620
rect 134380 56600 134620 56620
rect 134880 56600 135000 56620
rect 132000 56400 135000 56600
rect 132000 56380 132120 56400
rect 132380 56380 132620 56400
rect 132880 56380 133120 56400
rect 133380 56380 133620 56400
rect 133880 56380 134120 56400
rect 134380 56380 134620 56400
rect 134880 56380 135000 56400
rect 132000 56120 132100 56380
rect 132400 56120 132600 56380
rect 132900 56120 133100 56380
rect 133400 56120 133600 56380
rect 133900 56120 134100 56380
rect 134400 56120 134600 56380
rect 134900 56120 135000 56380
rect 132000 56100 132120 56120
rect 132380 56100 132620 56120
rect 132880 56100 133120 56120
rect 133380 56100 133620 56120
rect 133880 56100 134120 56120
rect 134380 56100 134620 56120
rect 134880 56100 135000 56120
rect 132000 55900 135000 56100
rect 132000 55880 132120 55900
rect 132380 55880 132620 55900
rect 132880 55880 133120 55900
rect 133380 55880 133620 55900
rect 133880 55880 134120 55900
rect 134380 55880 134620 55900
rect 134880 55880 135000 55900
rect 132000 55620 132100 55880
rect 132400 55620 132600 55880
rect 132900 55620 133100 55880
rect 133400 55620 133600 55880
rect 133900 55620 134100 55880
rect 134400 55620 134600 55880
rect 134900 55620 135000 55880
rect 132000 55600 132120 55620
rect 132380 55600 132620 55620
rect 132880 55600 133120 55620
rect 133380 55600 133620 55620
rect 133880 55600 134120 55620
rect 134380 55600 134620 55620
rect 134880 55600 135000 55620
rect 132000 55400 135000 55600
rect 132000 55380 132120 55400
rect 132380 55380 132620 55400
rect 132880 55380 133120 55400
rect 133380 55380 133620 55400
rect 133880 55380 134120 55400
rect 134380 55380 134620 55400
rect 134880 55380 135000 55400
rect 132000 55120 132100 55380
rect 132400 55120 132600 55380
rect 132900 55120 133100 55380
rect 133400 55120 133600 55380
rect 133900 55120 134100 55380
rect 134400 55120 134600 55380
rect 134900 55120 135000 55380
rect 132000 55100 132120 55120
rect 132380 55100 132620 55120
rect 132880 55100 133120 55120
rect 133380 55100 133620 55120
rect 133880 55100 134120 55120
rect 134380 55100 134620 55120
rect 134880 55100 135000 55120
rect 132000 54900 135000 55100
rect 132000 54880 132120 54900
rect 132380 54880 132620 54900
rect 132880 54880 133120 54900
rect 133380 54880 133620 54900
rect 133880 54880 134120 54900
rect 134380 54880 134620 54900
rect 134880 54880 135000 54900
rect 132000 54620 132100 54880
rect 132400 54620 132600 54880
rect 132900 54620 133100 54880
rect 133400 54620 133600 54880
rect 133900 54620 134100 54880
rect 134400 54620 134600 54880
rect 134900 54620 135000 54880
rect 132000 54600 132120 54620
rect 132380 54600 132620 54620
rect 132880 54600 133120 54620
rect 133380 54600 133620 54620
rect 133880 54600 134120 54620
rect 134380 54600 134620 54620
rect 134880 54600 135000 54620
rect 132000 54400 135000 54600
rect 132000 54380 132120 54400
rect 132380 54380 132620 54400
rect 132880 54380 133120 54400
rect 133380 54380 133620 54400
rect 133880 54380 134120 54400
rect 134380 54380 134620 54400
rect 134880 54380 135000 54400
rect 132000 54120 132100 54380
rect 132400 54120 132600 54380
rect 132900 54120 133100 54380
rect 133400 54120 133600 54380
rect 133900 54120 134100 54380
rect 134400 54120 134600 54380
rect 134900 54120 135000 54380
rect 132000 54100 132120 54120
rect 132380 54100 132620 54120
rect 132880 54100 133120 54120
rect 133380 54100 133620 54120
rect 133880 54100 134120 54120
rect 134380 54100 134620 54120
rect 134880 54100 135000 54120
rect 132000 53900 135000 54100
rect 132000 53880 132120 53900
rect 132380 53880 132620 53900
rect 132880 53880 133120 53900
rect 133380 53880 133620 53900
rect 133880 53880 134120 53900
rect 134380 53880 134620 53900
rect 134880 53880 135000 53900
rect 132000 53620 132100 53880
rect 132400 53620 132600 53880
rect 132900 53620 133100 53880
rect 133400 53620 133600 53880
rect 133900 53620 134100 53880
rect 134400 53620 134600 53880
rect 134900 53620 135000 53880
rect 132000 53600 132120 53620
rect 132380 53600 132620 53620
rect 132880 53600 133120 53620
rect 133380 53600 133620 53620
rect 133880 53600 134120 53620
rect 134380 53600 134620 53620
rect 134880 53600 135000 53620
rect 132000 53400 135000 53600
rect 132000 53380 132120 53400
rect 132380 53380 132620 53400
rect 132880 53380 133120 53400
rect 133380 53380 133620 53400
rect 133880 53380 134120 53400
rect 134380 53380 134620 53400
rect 134880 53380 135000 53400
rect 132000 53120 132100 53380
rect 132400 53120 132600 53380
rect 132900 53120 133100 53380
rect 133400 53120 133600 53380
rect 133900 53120 134100 53380
rect 134400 53120 134600 53380
rect 134900 53120 135000 53380
rect 132000 53100 132120 53120
rect 132380 53100 132620 53120
rect 132880 53100 133120 53120
rect 133380 53100 133620 53120
rect 133880 53100 134120 53120
rect 134380 53100 134620 53120
rect 134880 53100 135000 53120
rect 132000 52900 135000 53100
rect 132000 52880 132120 52900
rect 132380 52880 132620 52900
rect 132880 52880 133120 52900
rect 133380 52880 133620 52900
rect 133880 52880 134120 52900
rect 134380 52880 134620 52900
rect 134880 52880 135000 52900
rect 132000 52620 132100 52880
rect 132400 52620 132600 52880
rect 132900 52620 133100 52880
rect 133400 52620 133600 52880
rect 133900 52620 134100 52880
rect 134400 52620 134600 52880
rect 134900 52620 135000 52880
rect 132000 52600 132120 52620
rect 132380 52600 132620 52620
rect 132880 52600 133120 52620
rect 133380 52600 133620 52620
rect 133880 52600 134120 52620
rect 134380 52600 134620 52620
rect 134880 52600 135000 52620
rect 132000 52400 135000 52600
rect 132000 52380 132120 52400
rect 132380 52380 132620 52400
rect 132880 52380 133120 52400
rect 133380 52380 133620 52400
rect 133880 52380 134120 52400
rect 134380 52380 134620 52400
rect 134880 52380 135000 52400
rect 132000 52120 132100 52380
rect 132400 52120 132600 52380
rect 132900 52120 133100 52380
rect 133400 52120 133600 52380
rect 133900 52120 134100 52380
rect 134400 52120 134600 52380
rect 134900 52120 135000 52380
rect 132000 52100 132120 52120
rect 132380 52100 132620 52120
rect 132880 52100 133120 52120
rect 133380 52100 133620 52120
rect 133880 52100 134120 52120
rect 134380 52100 134620 52120
rect 134880 52100 135000 52120
rect 132000 51900 135000 52100
rect 132000 51880 132120 51900
rect 132380 51880 132620 51900
rect 132880 51880 133120 51900
rect 133380 51880 133620 51900
rect 133880 51880 134120 51900
rect 134380 51880 134620 51900
rect 134880 51880 135000 51900
rect 132000 51620 132100 51880
rect 132400 51620 132600 51880
rect 132900 51620 133100 51880
rect 133400 51620 133600 51880
rect 133900 51620 134100 51880
rect 134400 51620 134600 51880
rect 134900 51620 135000 51880
rect 132000 51600 132120 51620
rect 132380 51600 132620 51620
rect 132880 51600 133120 51620
rect 133380 51600 133620 51620
rect 133880 51600 134120 51620
rect 134380 51600 134620 51620
rect 134880 51600 135000 51620
rect 132000 51400 135000 51600
rect 132000 51380 132120 51400
rect 132380 51380 132620 51400
rect 132880 51380 133120 51400
rect 133380 51380 133620 51400
rect 133880 51380 134120 51400
rect 134380 51380 134620 51400
rect 134880 51380 135000 51400
rect 132000 51120 132100 51380
rect 132400 51120 132600 51380
rect 132900 51120 133100 51380
rect 133400 51120 133600 51380
rect 133900 51120 134100 51380
rect 134400 51120 134600 51380
rect 134900 51120 135000 51380
rect 132000 51100 132120 51120
rect 132380 51100 132620 51120
rect 132880 51100 133120 51120
rect 133380 51100 133620 51120
rect 133880 51100 134120 51120
rect 134380 51100 134620 51120
rect 134880 51100 135000 51120
rect 132000 50900 135000 51100
rect 132000 50880 132120 50900
rect 132380 50880 132620 50900
rect 132880 50880 133120 50900
rect 133380 50880 133620 50900
rect 133880 50880 134120 50900
rect 134380 50880 134620 50900
rect 134880 50880 135000 50900
rect 132000 50620 132100 50880
rect 132400 50620 132600 50880
rect 132900 50620 133100 50880
rect 133400 50620 133600 50880
rect 133900 50620 134100 50880
rect 134400 50620 134600 50880
rect 134900 50620 135000 50880
rect 132000 50600 132120 50620
rect 132380 50600 132620 50620
rect 132880 50600 133120 50620
rect 133380 50600 133620 50620
rect 133880 50600 134120 50620
rect 134380 50600 134620 50620
rect 134880 50600 135000 50620
rect 132000 50400 135000 50600
rect 132000 50380 132120 50400
rect 132380 50380 132620 50400
rect 132880 50380 133120 50400
rect 133380 50380 133620 50400
rect 133880 50380 134120 50400
rect 134380 50380 134620 50400
rect 134880 50380 135000 50400
rect 132000 50120 132100 50380
rect 132400 50120 132600 50380
rect 132900 50120 133100 50380
rect 133400 50120 133600 50380
rect 133900 50120 134100 50380
rect 134400 50120 134600 50380
rect 134900 50120 135000 50380
rect 132000 50100 132120 50120
rect 132380 50100 132620 50120
rect 132880 50100 133120 50120
rect 133380 50100 133620 50120
rect 133880 50100 134120 50120
rect 134380 50100 134620 50120
rect 134880 50100 135000 50120
rect 132000 49900 135000 50100
rect 132000 49880 132120 49900
rect 132380 49880 132620 49900
rect 132880 49880 133120 49900
rect 133380 49880 133620 49900
rect 133880 49880 134120 49900
rect 134380 49880 134620 49900
rect 134880 49880 135000 49900
rect 132000 49620 132100 49880
rect 132400 49620 132600 49880
rect 132900 49620 133100 49880
rect 133400 49620 133600 49880
rect 133900 49620 134100 49880
rect 134400 49620 134600 49880
rect 134900 49620 135000 49880
rect 132000 49600 132120 49620
rect 132380 49600 132620 49620
rect 132880 49600 133120 49620
rect 133380 49600 133620 49620
rect 133880 49600 134120 49620
rect 134380 49600 134620 49620
rect 134880 49600 135000 49620
rect 132000 49400 135000 49600
rect 132000 49380 132120 49400
rect 132380 49380 132620 49400
rect 132880 49380 133120 49400
rect 133380 49380 133620 49400
rect 133880 49380 134120 49400
rect 134380 49380 134620 49400
rect 134880 49380 135000 49400
rect 132000 49120 132100 49380
rect 132400 49120 132600 49380
rect 132900 49120 133100 49380
rect 133400 49120 133600 49380
rect 133900 49120 134100 49380
rect 134400 49120 134600 49380
rect 134900 49120 135000 49380
rect 132000 49100 132120 49120
rect 132380 49100 132620 49120
rect 132880 49100 133120 49120
rect 133380 49100 133620 49120
rect 133880 49100 134120 49120
rect 134380 49100 134620 49120
rect 134880 49100 135000 49120
rect 132000 48900 135000 49100
rect 132000 48880 132120 48900
rect 132380 48880 132620 48900
rect 132880 48880 133120 48900
rect 133380 48880 133620 48900
rect 133880 48880 134120 48900
rect 134380 48880 134620 48900
rect 134880 48880 135000 48900
rect 132000 48620 132100 48880
rect 132400 48620 132600 48880
rect 132900 48620 133100 48880
rect 133400 48620 133600 48880
rect 133900 48620 134100 48880
rect 134400 48620 134600 48880
rect 134900 48620 135000 48880
rect 132000 48600 132120 48620
rect 132380 48600 132620 48620
rect 132880 48600 133120 48620
rect 133380 48600 133620 48620
rect 133880 48600 134120 48620
rect 134380 48600 134620 48620
rect 134880 48600 135000 48620
rect 132000 48400 135000 48600
rect 132000 48380 132120 48400
rect 132380 48380 132620 48400
rect 132880 48380 133120 48400
rect 133380 48380 133620 48400
rect 133880 48380 134120 48400
rect 134380 48380 134620 48400
rect 134880 48380 135000 48400
rect 132000 48120 132100 48380
rect 132400 48120 132600 48380
rect 132900 48120 133100 48380
rect 133400 48120 133600 48380
rect 133900 48120 134100 48380
rect 134400 48120 134600 48380
rect 134900 48120 135000 48380
rect 132000 48100 132120 48120
rect 132380 48100 132620 48120
rect 132880 48100 133120 48120
rect 133380 48100 133620 48120
rect 133880 48100 134120 48120
rect 134380 48100 134620 48120
rect 134880 48100 135000 48120
rect 132000 47900 135000 48100
rect 132000 47880 132120 47900
rect 132380 47880 132620 47900
rect 132880 47880 133120 47900
rect 133380 47880 133620 47900
rect 133880 47880 134120 47900
rect 134380 47880 134620 47900
rect 134880 47880 135000 47900
rect 132000 47620 132100 47880
rect 132400 47620 132600 47880
rect 132900 47620 133100 47880
rect 133400 47620 133600 47880
rect 133900 47620 134100 47880
rect 134400 47620 134600 47880
rect 134900 47620 135000 47880
rect 132000 47600 132120 47620
rect 132380 47600 132620 47620
rect 132880 47600 133120 47620
rect 133380 47600 133620 47620
rect 133880 47600 134120 47620
rect 134380 47600 134620 47620
rect 134880 47600 135000 47620
rect 132000 47400 135000 47600
rect 132000 47380 132120 47400
rect 132380 47380 132620 47400
rect 132880 47380 133120 47400
rect 133380 47380 133620 47400
rect 133880 47380 134120 47400
rect 134380 47380 134620 47400
rect 134880 47380 135000 47400
rect 132000 47120 132100 47380
rect 132400 47120 132600 47380
rect 132900 47120 133100 47380
rect 133400 47120 133600 47380
rect 133900 47120 134100 47380
rect 134400 47120 134600 47380
rect 134900 47120 135000 47380
rect 132000 47100 132120 47120
rect 132380 47100 132620 47120
rect 132880 47100 133120 47120
rect 133380 47100 133620 47120
rect 133880 47100 134120 47120
rect 134380 47100 134620 47120
rect 134880 47100 135000 47120
rect 132000 46900 135000 47100
rect 132000 46880 132120 46900
rect 132380 46880 132620 46900
rect 132880 46880 133120 46900
rect 133380 46880 133620 46900
rect 133880 46880 134120 46900
rect 134380 46880 134620 46900
rect 134880 46880 135000 46900
rect 132000 46620 132100 46880
rect 132400 46620 132600 46880
rect 132900 46620 133100 46880
rect 133400 46620 133600 46880
rect 133900 46620 134100 46880
rect 134400 46620 134600 46880
rect 134900 46620 135000 46880
rect 132000 46600 132120 46620
rect 132380 46600 132620 46620
rect 132880 46600 133120 46620
rect 133380 46600 133620 46620
rect 133880 46600 134120 46620
rect 134380 46600 134620 46620
rect 134880 46600 135000 46620
rect 132000 46400 135000 46600
rect 132000 46380 132120 46400
rect 132380 46380 132620 46400
rect 132880 46380 133120 46400
rect 133380 46380 133620 46400
rect 133880 46380 134120 46400
rect 134380 46380 134620 46400
rect 134880 46380 135000 46400
rect 132000 46120 132100 46380
rect 132400 46120 132600 46380
rect 132900 46120 133100 46380
rect 133400 46120 133600 46380
rect 133900 46120 134100 46380
rect 134400 46120 134600 46380
rect 134900 46120 135000 46380
rect 132000 46100 132120 46120
rect 132380 46100 132620 46120
rect 132880 46100 133120 46120
rect 133380 46100 133620 46120
rect 133880 46100 134120 46120
rect 134380 46100 134620 46120
rect 134880 46100 135000 46120
rect 132000 45900 135000 46100
rect 132000 45880 132120 45900
rect 132380 45880 132620 45900
rect 132880 45880 133120 45900
rect 133380 45880 133620 45900
rect 133880 45880 134120 45900
rect 134380 45880 134620 45900
rect 134880 45880 135000 45900
rect 132000 45620 132100 45880
rect 132400 45620 132600 45880
rect 132900 45620 133100 45880
rect 133400 45620 133600 45880
rect 133900 45620 134100 45880
rect 134400 45620 134600 45880
rect 134900 45620 135000 45880
rect 132000 45600 132120 45620
rect 132380 45600 132620 45620
rect 132880 45600 133120 45620
rect 133380 45600 133620 45620
rect 133880 45600 134120 45620
rect 134380 45600 134620 45620
rect 134880 45600 135000 45620
rect 132000 45400 135000 45600
rect 132000 45380 132120 45400
rect 132380 45380 132620 45400
rect 132880 45380 133120 45400
rect 133380 45380 133620 45400
rect 133880 45380 134120 45400
rect 134380 45380 134620 45400
rect 134880 45380 135000 45400
rect 132000 45120 132100 45380
rect 132400 45120 132600 45380
rect 132900 45120 133100 45380
rect 133400 45120 133600 45380
rect 133900 45120 134100 45380
rect 134400 45120 134600 45380
rect 134900 45120 135000 45380
rect 132000 45100 132120 45120
rect 132380 45100 132620 45120
rect 132880 45100 133120 45120
rect 133380 45100 133620 45120
rect 133880 45100 134120 45120
rect 134380 45100 134620 45120
rect 134880 45100 135000 45120
rect 132000 44900 135000 45100
rect 132000 44880 132120 44900
rect 132380 44880 132620 44900
rect 132880 44880 133120 44900
rect 133380 44880 133620 44900
rect 133880 44880 134120 44900
rect 134380 44880 134620 44900
rect 134880 44880 135000 44900
rect 132000 44620 132100 44880
rect 132400 44620 132600 44880
rect 132900 44620 133100 44880
rect 133400 44620 133600 44880
rect 133900 44620 134100 44880
rect 134400 44620 134600 44880
rect 134900 44620 135000 44880
rect 132000 44600 132120 44620
rect 132380 44600 132620 44620
rect 132880 44600 133120 44620
rect 133380 44600 133620 44620
rect 133880 44600 134120 44620
rect 134380 44600 134620 44620
rect 134880 44600 135000 44620
rect 132000 44400 135000 44600
rect 132000 44380 132120 44400
rect 132380 44380 132620 44400
rect 132880 44380 133120 44400
rect 133380 44380 133620 44400
rect 133880 44380 134120 44400
rect 134380 44380 134620 44400
rect 134880 44380 135000 44400
rect 132000 44120 132100 44380
rect 132400 44120 132600 44380
rect 132900 44120 133100 44380
rect 133400 44120 133600 44380
rect 133900 44120 134100 44380
rect 134400 44120 134600 44380
rect 134900 44120 135000 44380
rect 132000 44100 132120 44120
rect 132380 44100 132620 44120
rect 132880 44100 133120 44120
rect 133380 44100 133620 44120
rect 133880 44100 134120 44120
rect 134380 44100 134620 44120
rect 134880 44100 135000 44120
rect 132000 43900 135000 44100
rect 132000 43880 132120 43900
rect 132380 43880 132620 43900
rect 132880 43880 133120 43900
rect 133380 43880 133620 43900
rect 133880 43880 134120 43900
rect 134380 43880 134620 43900
rect 134880 43880 135000 43900
rect 132000 43620 132100 43880
rect 132400 43620 132600 43880
rect 132900 43620 133100 43880
rect 133400 43620 133600 43880
rect 133900 43620 134100 43880
rect 134400 43620 134600 43880
rect 134900 43620 135000 43880
rect 132000 43600 132120 43620
rect 132380 43600 132620 43620
rect 132880 43600 133120 43620
rect 133380 43600 133620 43620
rect 133880 43600 134120 43620
rect 134380 43600 134620 43620
rect 134880 43600 135000 43620
rect 132000 43400 135000 43600
rect 132000 43380 132120 43400
rect 132380 43380 132620 43400
rect 132880 43380 133120 43400
rect 133380 43380 133620 43400
rect 133880 43380 134120 43400
rect 134380 43380 134620 43400
rect 134880 43380 135000 43400
rect 132000 43120 132100 43380
rect 132400 43120 132600 43380
rect 132900 43120 133100 43380
rect 133400 43120 133600 43380
rect 133900 43120 134100 43380
rect 134400 43120 134600 43380
rect 134900 43120 135000 43380
rect 132000 43100 132120 43120
rect 132380 43100 132620 43120
rect 132880 43100 133120 43120
rect 133380 43100 133620 43120
rect 133880 43100 134120 43120
rect 134380 43100 134620 43120
rect 134880 43100 135000 43120
rect 132000 42900 135000 43100
rect 132000 42880 132120 42900
rect 132380 42880 132620 42900
rect 132880 42880 133120 42900
rect 133380 42880 133620 42900
rect 133880 42880 134120 42900
rect 134380 42880 134620 42900
rect 134880 42880 135000 42900
rect 132000 42620 132100 42880
rect 132400 42620 132600 42880
rect 132900 42620 133100 42880
rect 133400 42620 133600 42880
rect 133900 42620 134100 42880
rect 134400 42620 134600 42880
rect 134900 42620 135000 42880
rect 132000 42600 132120 42620
rect 132380 42600 132620 42620
rect 132880 42600 133120 42620
rect 133380 42600 133620 42620
rect 133880 42600 134120 42620
rect 134380 42600 134620 42620
rect 134880 42600 135000 42620
rect 132000 42400 135000 42600
rect 132000 42380 132120 42400
rect 132380 42380 132620 42400
rect 132880 42380 133120 42400
rect 133380 42380 133620 42400
rect 133880 42380 134120 42400
rect 134380 42380 134620 42400
rect 134880 42380 135000 42400
rect 132000 42120 132100 42380
rect 132400 42120 132600 42380
rect 132900 42120 133100 42380
rect 133400 42120 133600 42380
rect 133900 42120 134100 42380
rect 134400 42120 134600 42380
rect 134900 42120 135000 42380
rect 132000 42100 132120 42120
rect 132380 42100 132620 42120
rect 132880 42100 133120 42120
rect 133380 42100 133620 42120
rect 133880 42100 134120 42120
rect 134380 42100 134620 42120
rect 134880 42100 135000 42120
rect 132000 41900 135000 42100
rect 132000 41880 132120 41900
rect 132380 41880 132620 41900
rect 132880 41880 133120 41900
rect 133380 41880 133620 41900
rect 133880 41880 134120 41900
rect 134380 41880 134620 41900
rect 134880 41880 135000 41900
rect 132000 41620 132100 41880
rect 132400 41620 132600 41880
rect 132900 41620 133100 41880
rect 133400 41620 133600 41880
rect 133900 41620 134100 41880
rect 134400 41620 134600 41880
rect 134900 41620 135000 41880
rect 132000 41600 132120 41620
rect 132380 41600 132620 41620
rect 132880 41600 133120 41620
rect 133380 41600 133620 41620
rect 133880 41600 134120 41620
rect 134380 41600 134620 41620
rect 134880 41600 135000 41620
rect 132000 41400 135000 41600
rect 132000 41380 132120 41400
rect 132380 41380 132620 41400
rect 132880 41380 133120 41400
rect 133380 41380 133620 41400
rect 133880 41380 134120 41400
rect 134380 41380 134620 41400
rect 134880 41380 135000 41400
rect 132000 41120 132100 41380
rect 132400 41120 132600 41380
rect 132900 41120 133100 41380
rect 133400 41120 133600 41380
rect 133900 41120 134100 41380
rect 134400 41120 134600 41380
rect 134900 41120 135000 41380
rect 132000 41100 132120 41120
rect 132380 41100 132620 41120
rect 132880 41100 133120 41120
rect 133380 41100 133620 41120
rect 133880 41100 134120 41120
rect 134380 41100 134620 41120
rect 134880 41100 135000 41120
rect 132000 40900 135000 41100
rect 132000 40880 132120 40900
rect 132380 40880 132620 40900
rect 132880 40880 133120 40900
rect 133380 40880 133620 40900
rect 133880 40880 134120 40900
rect 134380 40880 134620 40900
rect 134880 40880 135000 40900
rect 132000 40620 132100 40880
rect 132400 40620 132600 40880
rect 132900 40620 133100 40880
rect 133400 40620 133600 40880
rect 133900 40620 134100 40880
rect 134400 40620 134600 40880
rect 134900 40620 135000 40880
rect 132000 40600 132120 40620
rect 132380 40600 132620 40620
rect 132880 40600 133120 40620
rect 133380 40600 133620 40620
rect 133880 40600 134120 40620
rect 134380 40600 134620 40620
rect 134880 40600 135000 40620
rect 132000 40400 135000 40600
rect 132000 40380 132120 40400
rect 132380 40380 132620 40400
rect 132880 40380 133120 40400
rect 133380 40380 133620 40400
rect 133880 40380 134120 40400
rect 134380 40380 134620 40400
rect 134880 40380 135000 40400
rect 132000 40120 132100 40380
rect 132400 40120 132600 40380
rect 132900 40120 133100 40380
rect 133400 40120 133600 40380
rect 133900 40120 134100 40380
rect 134400 40120 134600 40380
rect 134900 40120 135000 40380
rect 132000 40100 132120 40120
rect 132380 40100 132620 40120
rect 132880 40100 133120 40120
rect 133380 40100 133620 40120
rect 133880 40100 134120 40120
rect 134380 40100 134620 40120
rect 134880 40100 135000 40120
rect 132000 39900 135000 40100
rect 132000 39880 132120 39900
rect 132380 39880 132620 39900
rect 132880 39880 133120 39900
rect 133380 39880 133620 39900
rect 133880 39880 134120 39900
rect 134380 39880 134620 39900
rect 134880 39880 135000 39900
rect 132000 39620 132100 39880
rect 132400 39620 132600 39880
rect 132900 39620 133100 39880
rect 133400 39620 133600 39880
rect 133900 39620 134100 39880
rect 134400 39620 134600 39880
rect 134900 39620 135000 39880
rect 132000 39600 132120 39620
rect 132380 39600 132620 39620
rect 132880 39600 133120 39620
rect 133380 39600 133620 39620
rect 133880 39600 134120 39620
rect 134380 39600 134620 39620
rect 134880 39600 135000 39620
rect 132000 39400 135000 39600
rect 132000 39380 132120 39400
rect 132380 39380 132620 39400
rect 132880 39380 133120 39400
rect 133380 39380 133620 39400
rect 133880 39380 134120 39400
rect 134380 39380 134620 39400
rect 134880 39380 135000 39400
rect 132000 39120 132100 39380
rect 132400 39120 132600 39380
rect 132900 39120 133100 39380
rect 133400 39120 133600 39380
rect 133900 39120 134100 39380
rect 134400 39120 134600 39380
rect 134900 39120 135000 39380
rect 132000 39100 132120 39120
rect 132380 39100 132620 39120
rect 132880 39100 133120 39120
rect 133380 39100 133620 39120
rect 133880 39100 134120 39120
rect 134380 39100 134620 39120
rect 134880 39100 135000 39120
rect 132000 39000 135000 39100
rect 204000 63980 208000 64000
rect 204000 63910 204150 63980
rect 204350 63910 204650 63980
rect 204850 63910 205150 63980
rect 205350 63910 205650 63980
rect 205850 63910 206150 63980
rect 206350 63910 206650 63980
rect 206850 63910 207150 63980
rect 207350 63910 207650 63980
rect 207850 63910 208000 63980
rect 204000 63900 208000 63910
rect 204000 63880 204120 63900
rect 204380 63880 204620 63900
rect 204880 63880 205120 63900
rect 205380 63880 205620 63900
rect 205880 63880 206120 63900
rect 206380 63880 206620 63900
rect 206880 63880 207120 63900
rect 207380 63880 207620 63900
rect 207880 63880 208000 63900
rect 204000 63850 204100 63880
rect 204000 63650 204020 63850
rect 204090 63650 204100 63850
rect 204000 63620 204100 63650
rect 204400 63850 204600 63880
rect 204400 63650 204410 63850
rect 204480 63650 204520 63850
rect 204590 63650 204600 63850
rect 204400 63620 204600 63650
rect 204900 63850 205100 63880
rect 204900 63650 204910 63850
rect 204980 63650 205020 63850
rect 205090 63650 205100 63850
rect 204900 63620 205100 63650
rect 205400 63850 205600 63880
rect 205400 63650 205410 63850
rect 205480 63650 205520 63850
rect 205590 63650 205600 63850
rect 205400 63620 205600 63650
rect 205900 63850 206100 63880
rect 205900 63650 205910 63850
rect 205980 63650 206020 63850
rect 206090 63650 206100 63850
rect 205900 63620 206100 63650
rect 206400 63850 206600 63880
rect 206400 63650 206410 63850
rect 206480 63650 206520 63850
rect 206590 63650 206600 63850
rect 206400 63620 206600 63650
rect 206900 63850 207100 63880
rect 206900 63650 206910 63850
rect 206980 63650 207020 63850
rect 207090 63650 207100 63850
rect 206900 63620 207100 63650
rect 207400 63850 207600 63880
rect 207400 63650 207410 63850
rect 207480 63650 207520 63850
rect 207590 63650 207600 63850
rect 207400 63620 207600 63650
rect 207900 63850 208000 63880
rect 207900 63650 207910 63850
rect 207980 63650 208000 63850
rect 207900 63620 208000 63650
rect 204000 63600 204120 63620
rect 204380 63600 204620 63620
rect 204880 63600 205120 63620
rect 205380 63600 205620 63620
rect 205880 63600 206120 63620
rect 206380 63600 206620 63620
rect 206880 63600 207120 63620
rect 207380 63600 207620 63620
rect 207880 63600 208000 63620
rect 204000 63590 208000 63600
rect 204000 63520 204150 63590
rect 204350 63520 204650 63590
rect 204850 63520 205150 63590
rect 205350 63520 205650 63590
rect 205850 63520 206150 63590
rect 206350 63520 206650 63590
rect 206850 63520 207150 63590
rect 207350 63520 207650 63590
rect 207850 63520 208000 63590
rect 204000 63480 208000 63520
rect 204000 63410 204150 63480
rect 204350 63410 204650 63480
rect 204850 63410 205150 63480
rect 205350 63410 205650 63480
rect 205850 63410 206150 63480
rect 206350 63410 206650 63480
rect 206850 63410 207150 63480
rect 207350 63410 207650 63480
rect 207850 63410 208000 63480
rect 204000 63400 208000 63410
rect 204000 63380 204120 63400
rect 204380 63380 204620 63400
rect 204880 63380 205120 63400
rect 205380 63380 205620 63400
rect 205880 63380 206120 63400
rect 206380 63380 206620 63400
rect 206880 63380 207120 63400
rect 207380 63380 207620 63400
rect 207880 63380 208000 63400
rect 204000 63350 204100 63380
rect 204000 63150 204020 63350
rect 204090 63150 204100 63350
rect 204000 63120 204100 63150
rect 204400 63350 204600 63380
rect 204400 63150 204410 63350
rect 204480 63150 204520 63350
rect 204590 63150 204600 63350
rect 204400 63120 204600 63150
rect 204900 63350 205100 63380
rect 204900 63150 204910 63350
rect 204980 63150 205020 63350
rect 205090 63150 205100 63350
rect 204900 63120 205100 63150
rect 205400 63350 205600 63380
rect 205400 63150 205410 63350
rect 205480 63150 205520 63350
rect 205590 63150 205600 63350
rect 205400 63120 205600 63150
rect 205900 63350 206100 63380
rect 205900 63150 205910 63350
rect 205980 63150 206020 63350
rect 206090 63150 206100 63350
rect 205900 63120 206100 63150
rect 206400 63350 206600 63380
rect 206400 63150 206410 63350
rect 206480 63150 206520 63350
rect 206590 63150 206600 63350
rect 206400 63120 206600 63150
rect 206900 63350 207100 63380
rect 206900 63150 206910 63350
rect 206980 63150 207020 63350
rect 207090 63150 207100 63350
rect 206900 63120 207100 63150
rect 207400 63350 207600 63380
rect 207400 63150 207410 63350
rect 207480 63150 207520 63350
rect 207590 63150 207600 63350
rect 207400 63120 207600 63150
rect 207900 63350 208000 63380
rect 207900 63150 207910 63350
rect 207980 63150 208000 63350
rect 207900 63120 208000 63150
rect 204000 63100 204120 63120
rect 204380 63100 204620 63120
rect 204880 63100 205120 63120
rect 205380 63100 205620 63120
rect 205880 63100 206120 63120
rect 206380 63100 206620 63120
rect 206880 63100 207120 63120
rect 207380 63100 207620 63120
rect 207880 63100 208000 63120
rect 204000 63090 208000 63100
rect 204000 63020 204150 63090
rect 204350 63020 204650 63090
rect 204850 63020 205150 63090
rect 205350 63020 205650 63090
rect 205850 63020 206150 63090
rect 206350 63020 206650 63090
rect 206850 63020 207150 63090
rect 207350 63020 207650 63090
rect 207850 63020 208000 63090
rect 204000 62980 208000 63020
rect 204000 62910 204150 62980
rect 204350 62910 204650 62980
rect 204850 62910 205150 62980
rect 205350 62910 205650 62980
rect 205850 62910 206150 62980
rect 206350 62910 206650 62980
rect 206850 62910 207150 62980
rect 207350 62910 207650 62980
rect 207850 62910 208000 62980
rect 204000 62900 208000 62910
rect 204000 62880 204120 62900
rect 204380 62880 204620 62900
rect 204880 62880 205120 62900
rect 205380 62880 205620 62900
rect 205880 62880 206120 62900
rect 206380 62880 206620 62900
rect 206880 62880 207120 62900
rect 207380 62880 207620 62900
rect 207880 62880 208000 62900
rect 204000 62850 204100 62880
rect 204000 62650 204020 62850
rect 204090 62650 204100 62850
rect 204000 62620 204100 62650
rect 204400 62850 204600 62880
rect 204400 62650 204410 62850
rect 204480 62650 204520 62850
rect 204590 62650 204600 62850
rect 204400 62620 204600 62650
rect 204900 62850 205100 62880
rect 204900 62650 204910 62850
rect 204980 62650 205020 62850
rect 205090 62650 205100 62850
rect 204900 62620 205100 62650
rect 205400 62850 205600 62880
rect 205400 62650 205410 62850
rect 205480 62650 205520 62850
rect 205590 62650 205600 62850
rect 205400 62620 205600 62650
rect 205900 62850 206100 62880
rect 205900 62650 205910 62850
rect 205980 62650 206020 62850
rect 206090 62650 206100 62850
rect 205900 62620 206100 62650
rect 206400 62850 206600 62880
rect 206400 62650 206410 62850
rect 206480 62650 206520 62850
rect 206590 62650 206600 62850
rect 206400 62620 206600 62650
rect 206900 62850 207100 62880
rect 206900 62650 206910 62850
rect 206980 62650 207020 62850
rect 207090 62650 207100 62850
rect 206900 62620 207100 62650
rect 207400 62850 207600 62880
rect 207400 62650 207410 62850
rect 207480 62650 207520 62850
rect 207590 62650 207600 62850
rect 207400 62620 207600 62650
rect 207900 62850 208000 62880
rect 207900 62650 207910 62850
rect 207980 62650 208000 62850
rect 207900 62620 208000 62650
rect 204000 62600 204120 62620
rect 204380 62600 204620 62620
rect 204880 62600 205120 62620
rect 205380 62600 205620 62620
rect 205880 62600 206120 62620
rect 206380 62600 206620 62620
rect 206880 62600 207120 62620
rect 207380 62600 207620 62620
rect 207880 62600 208000 62620
rect 204000 62590 208000 62600
rect 204000 62520 204150 62590
rect 204350 62520 204650 62590
rect 204850 62520 205150 62590
rect 205350 62520 205650 62590
rect 205850 62520 206150 62590
rect 206350 62520 206650 62590
rect 206850 62520 207150 62590
rect 207350 62520 207650 62590
rect 207850 62520 208000 62590
rect 204000 62480 208000 62520
rect 204000 62410 204150 62480
rect 204350 62410 204650 62480
rect 204850 62410 205150 62480
rect 205350 62410 205650 62480
rect 205850 62410 206150 62480
rect 206350 62410 206650 62480
rect 206850 62410 207150 62480
rect 207350 62410 207650 62480
rect 207850 62410 208000 62480
rect 204000 62400 208000 62410
rect 204000 62380 204120 62400
rect 204380 62380 204620 62400
rect 204880 62380 205120 62400
rect 205380 62380 205620 62400
rect 205880 62380 206120 62400
rect 206380 62380 206620 62400
rect 206880 62380 207120 62400
rect 207380 62380 207620 62400
rect 207880 62380 208000 62400
rect 204000 62350 204100 62380
rect 204000 62150 204020 62350
rect 204090 62150 204100 62350
rect 204000 62120 204100 62150
rect 204400 62350 204600 62380
rect 204400 62150 204410 62350
rect 204480 62150 204520 62350
rect 204590 62150 204600 62350
rect 204400 62120 204600 62150
rect 204900 62350 205100 62380
rect 204900 62150 204910 62350
rect 204980 62150 205020 62350
rect 205090 62150 205100 62350
rect 204900 62120 205100 62150
rect 205400 62350 205600 62380
rect 205400 62150 205410 62350
rect 205480 62150 205520 62350
rect 205590 62150 205600 62350
rect 205400 62120 205600 62150
rect 205900 62350 206100 62380
rect 205900 62150 205910 62350
rect 205980 62150 206020 62350
rect 206090 62150 206100 62350
rect 205900 62120 206100 62150
rect 206400 62350 206600 62380
rect 206400 62150 206410 62350
rect 206480 62150 206520 62350
rect 206590 62150 206600 62350
rect 206400 62120 206600 62150
rect 206900 62350 207100 62380
rect 206900 62150 206910 62350
rect 206980 62150 207020 62350
rect 207090 62150 207100 62350
rect 206900 62120 207100 62150
rect 207400 62350 207600 62380
rect 207400 62150 207410 62350
rect 207480 62150 207520 62350
rect 207590 62150 207600 62350
rect 207400 62120 207600 62150
rect 207900 62350 208000 62380
rect 207900 62150 207910 62350
rect 207980 62150 208000 62350
rect 207900 62120 208000 62150
rect 204000 62100 204120 62120
rect 204380 62100 204620 62120
rect 204880 62100 205120 62120
rect 205380 62100 205620 62120
rect 205880 62100 206120 62120
rect 206380 62100 206620 62120
rect 206880 62100 207120 62120
rect 207380 62100 207620 62120
rect 207880 62100 208000 62120
rect 204000 62090 208000 62100
rect 204000 62020 204150 62090
rect 204350 62020 204650 62090
rect 204850 62020 205150 62090
rect 205350 62020 205650 62090
rect 205850 62020 206150 62090
rect 206350 62020 206650 62090
rect 206850 62020 207150 62090
rect 207350 62020 207650 62090
rect 207850 62020 208000 62090
rect 204000 61980 208000 62020
rect 204000 61910 204150 61980
rect 204350 61910 204650 61980
rect 204850 61910 205150 61980
rect 205350 61910 205650 61980
rect 205850 61910 206150 61980
rect 206350 61910 206650 61980
rect 206850 61910 207150 61980
rect 207350 61910 207650 61980
rect 207850 61910 208000 61980
rect 204000 61900 208000 61910
rect 204000 61880 204120 61900
rect 204380 61880 204620 61900
rect 204880 61880 205120 61900
rect 205380 61880 205620 61900
rect 205880 61880 206120 61900
rect 206380 61880 206620 61900
rect 206880 61880 207120 61900
rect 207380 61880 207620 61900
rect 207880 61880 208000 61900
rect 204000 61850 204100 61880
rect 204000 61650 204020 61850
rect 204090 61650 204100 61850
rect 204000 61620 204100 61650
rect 204400 61850 204600 61880
rect 204400 61650 204410 61850
rect 204480 61650 204520 61850
rect 204590 61650 204600 61850
rect 204400 61620 204600 61650
rect 204900 61850 205100 61880
rect 204900 61650 204910 61850
rect 204980 61650 205020 61850
rect 205090 61650 205100 61850
rect 204900 61620 205100 61650
rect 205400 61850 205600 61880
rect 205400 61650 205410 61850
rect 205480 61650 205520 61850
rect 205590 61650 205600 61850
rect 205400 61620 205600 61650
rect 205900 61850 206100 61880
rect 205900 61650 205910 61850
rect 205980 61650 206020 61850
rect 206090 61650 206100 61850
rect 205900 61620 206100 61650
rect 206400 61850 206600 61880
rect 206400 61650 206410 61850
rect 206480 61650 206520 61850
rect 206590 61650 206600 61850
rect 206400 61620 206600 61650
rect 206900 61850 207100 61880
rect 206900 61650 206910 61850
rect 206980 61650 207020 61850
rect 207090 61650 207100 61850
rect 206900 61620 207100 61650
rect 207400 61850 207600 61880
rect 207400 61650 207410 61850
rect 207480 61650 207520 61850
rect 207590 61650 207600 61850
rect 207400 61620 207600 61650
rect 207900 61850 208000 61880
rect 207900 61650 207910 61850
rect 207980 61650 208000 61850
rect 207900 61620 208000 61650
rect 204000 61600 204120 61620
rect 204380 61600 204620 61620
rect 204880 61600 205120 61620
rect 205380 61600 205620 61620
rect 205880 61600 206120 61620
rect 206380 61600 206620 61620
rect 206880 61600 207120 61620
rect 207380 61600 207620 61620
rect 207880 61600 208000 61620
rect 204000 61590 208000 61600
rect 204000 61520 204150 61590
rect 204350 61520 204650 61590
rect 204850 61520 205150 61590
rect 205350 61520 205650 61590
rect 205850 61520 206150 61590
rect 206350 61520 206650 61590
rect 206850 61520 207150 61590
rect 207350 61520 207650 61590
rect 207850 61520 208000 61590
rect 204000 61480 208000 61520
rect 204000 61410 204150 61480
rect 204350 61410 204650 61480
rect 204850 61410 205150 61480
rect 205350 61410 205650 61480
rect 205850 61410 206150 61480
rect 206350 61410 206650 61480
rect 206850 61410 207150 61480
rect 207350 61410 207650 61480
rect 207850 61410 208000 61480
rect 204000 61400 208000 61410
rect 204000 61380 204120 61400
rect 204380 61380 204620 61400
rect 204880 61380 205120 61400
rect 205380 61380 205620 61400
rect 205880 61380 206120 61400
rect 206380 61380 206620 61400
rect 206880 61380 207120 61400
rect 207380 61380 207620 61400
rect 207880 61380 208000 61400
rect 204000 61350 204100 61380
rect 204000 61150 204020 61350
rect 204090 61150 204100 61350
rect 204000 61120 204100 61150
rect 204400 61350 204600 61380
rect 204400 61150 204410 61350
rect 204480 61150 204520 61350
rect 204590 61150 204600 61350
rect 204400 61120 204600 61150
rect 204900 61350 205100 61380
rect 204900 61150 204910 61350
rect 204980 61150 205020 61350
rect 205090 61150 205100 61350
rect 204900 61120 205100 61150
rect 205400 61350 205600 61380
rect 205400 61150 205410 61350
rect 205480 61150 205520 61350
rect 205590 61150 205600 61350
rect 205400 61120 205600 61150
rect 205900 61350 206100 61380
rect 205900 61150 205910 61350
rect 205980 61150 206020 61350
rect 206090 61150 206100 61350
rect 205900 61120 206100 61150
rect 206400 61350 206600 61380
rect 206400 61150 206410 61350
rect 206480 61150 206520 61350
rect 206590 61150 206600 61350
rect 206400 61120 206600 61150
rect 206900 61350 207100 61380
rect 206900 61150 206910 61350
rect 206980 61150 207020 61350
rect 207090 61150 207100 61350
rect 206900 61120 207100 61150
rect 207400 61350 207600 61380
rect 207400 61150 207410 61350
rect 207480 61150 207520 61350
rect 207590 61150 207600 61350
rect 207400 61120 207600 61150
rect 207900 61350 208000 61380
rect 207900 61150 207910 61350
rect 207980 61150 208000 61350
rect 207900 61120 208000 61150
rect 204000 61100 204120 61120
rect 204380 61100 204620 61120
rect 204880 61100 205120 61120
rect 205380 61100 205620 61120
rect 205880 61100 206120 61120
rect 206380 61100 206620 61120
rect 206880 61100 207120 61120
rect 207380 61100 207620 61120
rect 207880 61100 208000 61120
rect 204000 61090 208000 61100
rect 204000 61020 204150 61090
rect 204350 61020 204650 61090
rect 204850 61020 205150 61090
rect 205350 61020 205650 61090
rect 205850 61020 206150 61090
rect 206350 61020 206650 61090
rect 206850 61020 207150 61090
rect 207350 61020 207650 61090
rect 207850 61020 208000 61090
rect 204000 60980 208000 61020
rect 204000 60910 204150 60980
rect 204350 60910 204650 60980
rect 204850 60910 205150 60980
rect 205350 60910 205650 60980
rect 205850 60910 206150 60980
rect 206350 60910 206650 60980
rect 206850 60910 207150 60980
rect 207350 60910 207650 60980
rect 207850 60910 208000 60980
rect 204000 60900 208000 60910
rect 204000 60880 204120 60900
rect 204380 60880 204620 60900
rect 204880 60880 205120 60900
rect 205380 60880 205620 60900
rect 205880 60880 206120 60900
rect 206380 60880 206620 60900
rect 206880 60880 207120 60900
rect 207380 60880 207620 60900
rect 207880 60880 208000 60900
rect 204000 60850 204100 60880
rect 204000 60650 204020 60850
rect 204090 60650 204100 60850
rect 204000 60620 204100 60650
rect 204400 60850 204600 60880
rect 204400 60650 204410 60850
rect 204480 60650 204520 60850
rect 204590 60650 204600 60850
rect 204400 60620 204600 60650
rect 204900 60850 205100 60880
rect 204900 60650 204910 60850
rect 204980 60650 205020 60850
rect 205090 60650 205100 60850
rect 204900 60620 205100 60650
rect 205400 60850 205600 60880
rect 205400 60650 205410 60850
rect 205480 60650 205520 60850
rect 205590 60650 205600 60850
rect 205400 60620 205600 60650
rect 205900 60850 206100 60880
rect 205900 60650 205910 60850
rect 205980 60650 206020 60850
rect 206090 60650 206100 60850
rect 205900 60620 206100 60650
rect 206400 60850 206600 60880
rect 206400 60650 206410 60850
rect 206480 60650 206520 60850
rect 206590 60650 206600 60850
rect 206400 60620 206600 60650
rect 206900 60850 207100 60880
rect 206900 60650 206910 60850
rect 206980 60650 207020 60850
rect 207090 60650 207100 60850
rect 206900 60620 207100 60650
rect 207400 60850 207600 60880
rect 207400 60650 207410 60850
rect 207480 60650 207520 60850
rect 207590 60650 207600 60850
rect 207400 60620 207600 60650
rect 207900 60850 208000 60880
rect 207900 60650 207910 60850
rect 207980 60650 208000 60850
rect 207900 60620 208000 60650
rect 204000 60600 204120 60620
rect 204380 60600 204620 60620
rect 204880 60600 205120 60620
rect 205380 60600 205620 60620
rect 205880 60600 206120 60620
rect 206380 60600 206620 60620
rect 206880 60600 207120 60620
rect 207380 60600 207620 60620
rect 207880 60600 208000 60620
rect 204000 60590 208000 60600
rect 204000 60520 204150 60590
rect 204350 60520 204650 60590
rect 204850 60520 205150 60590
rect 205350 60520 205650 60590
rect 205850 60520 206150 60590
rect 206350 60520 206650 60590
rect 206850 60520 207150 60590
rect 207350 60520 207650 60590
rect 207850 60520 208000 60590
rect 204000 60480 208000 60520
rect 204000 60410 204150 60480
rect 204350 60410 204650 60480
rect 204850 60410 205150 60480
rect 205350 60410 205650 60480
rect 205850 60410 206150 60480
rect 206350 60410 206650 60480
rect 206850 60410 207150 60480
rect 207350 60410 207650 60480
rect 207850 60410 208000 60480
rect 204000 60400 208000 60410
rect 204000 60380 204120 60400
rect 204380 60380 204620 60400
rect 204880 60380 205120 60400
rect 205380 60380 205620 60400
rect 205880 60380 206120 60400
rect 206380 60380 206620 60400
rect 206880 60380 207120 60400
rect 207380 60380 207620 60400
rect 207880 60380 208000 60400
rect 204000 60350 204100 60380
rect 204000 60150 204020 60350
rect 204090 60150 204100 60350
rect 204000 60120 204100 60150
rect 204400 60350 204600 60380
rect 204400 60150 204410 60350
rect 204480 60150 204520 60350
rect 204590 60150 204600 60350
rect 204400 60120 204600 60150
rect 204900 60350 205100 60380
rect 204900 60150 204910 60350
rect 204980 60150 205020 60350
rect 205090 60150 205100 60350
rect 204900 60120 205100 60150
rect 205400 60350 205600 60380
rect 205400 60150 205410 60350
rect 205480 60150 205520 60350
rect 205590 60150 205600 60350
rect 205400 60120 205600 60150
rect 205900 60350 206100 60380
rect 205900 60150 205910 60350
rect 205980 60150 206020 60350
rect 206090 60150 206100 60350
rect 205900 60120 206100 60150
rect 206400 60350 206600 60380
rect 206400 60150 206410 60350
rect 206480 60150 206520 60350
rect 206590 60150 206600 60350
rect 206400 60120 206600 60150
rect 206900 60350 207100 60380
rect 206900 60150 206910 60350
rect 206980 60150 207020 60350
rect 207090 60150 207100 60350
rect 206900 60120 207100 60150
rect 207400 60350 207600 60380
rect 207400 60150 207410 60350
rect 207480 60150 207520 60350
rect 207590 60150 207600 60350
rect 207400 60120 207600 60150
rect 207900 60350 208000 60380
rect 207900 60150 207910 60350
rect 207980 60150 208000 60350
rect 207900 60120 208000 60150
rect 204000 60100 204120 60120
rect 204380 60100 204620 60120
rect 204880 60100 205120 60120
rect 205380 60100 205620 60120
rect 205880 60100 206120 60120
rect 206380 60100 206620 60120
rect 206880 60100 207120 60120
rect 207380 60100 207620 60120
rect 207880 60100 208000 60120
rect 204000 60090 208000 60100
rect 204000 60020 204150 60090
rect 204350 60020 204650 60090
rect 204850 60020 205150 60090
rect 205350 60020 205650 60090
rect 205850 60020 206150 60090
rect 206350 60020 206650 60090
rect 206850 60020 207150 60090
rect 207350 60020 207650 60090
rect 207850 60020 208000 60090
rect 204000 59980 208000 60020
rect 204000 59910 204150 59980
rect 204350 59910 204650 59980
rect 204850 59910 205150 59980
rect 205350 59910 205650 59980
rect 205850 59910 206150 59980
rect 206350 59910 206650 59980
rect 206850 59910 207150 59980
rect 207350 59910 207650 59980
rect 207850 59910 208000 59980
rect 204000 59900 208000 59910
rect 204000 59880 204120 59900
rect 204380 59880 204620 59900
rect 204880 59880 205120 59900
rect 205380 59880 205620 59900
rect 205880 59880 206120 59900
rect 206380 59880 206620 59900
rect 206880 59880 207120 59900
rect 207380 59880 207620 59900
rect 207880 59880 208000 59900
rect 204000 59850 204100 59880
rect 204000 59650 204020 59850
rect 204090 59650 204100 59850
rect 204000 59620 204100 59650
rect 204400 59850 204600 59880
rect 204400 59650 204410 59850
rect 204480 59650 204520 59850
rect 204590 59650 204600 59850
rect 204400 59620 204600 59650
rect 204900 59850 205100 59880
rect 204900 59650 204910 59850
rect 204980 59650 205020 59850
rect 205090 59650 205100 59850
rect 204900 59620 205100 59650
rect 205400 59850 205600 59880
rect 205400 59650 205410 59850
rect 205480 59650 205520 59850
rect 205590 59650 205600 59850
rect 205400 59620 205600 59650
rect 205900 59850 206100 59880
rect 205900 59650 205910 59850
rect 205980 59650 206020 59850
rect 206090 59650 206100 59850
rect 205900 59620 206100 59650
rect 206400 59850 206600 59880
rect 206400 59650 206410 59850
rect 206480 59650 206520 59850
rect 206590 59650 206600 59850
rect 206400 59620 206600 59650
rect 206900 59850 207100 59880
rect 206900 59650 206910 59850
rect 206980 59650 207020 59850
rect 207090 59650 207100 59850
rect 206900 59620 207100 59650
rect 207400 59850 207600 59880
rect 207400 59650 207410 59850
rect 207480 59650 207520 59850
rect 207590 59650 207600 59850
rect 207400 59620 207600 59650
rect 207900 59850 208000 59880
rect 207900 59650 207910 59850
rect 207980 59650 208000 59850
rect 207900 59620 208000 59650
rect 204000 59600 204120 59620
rect 204380 59600 204620 59620
rect 204880 59600 205120 59620
rect 205380 59600 205620 59620
rect 205880 59600 206120 59620
rect 206380 59600 206620 59620
rect 206880 59600 207120 59620
rect 207380 59600 207620 59620
rect 207880 59600 208000 59620
rect 204000 59590 208000 59600
rect 204000 59520 204150 59590
rect 204350 59520 204650 59590
rect 204850 59520 205150 59590
rect 205350 59520 205650 59590
rect 205850 59520 206150 59590
rect 206350 59520 206650 59590
rect 206850 59520 207150 59590
rect 207350 59520 207650 59590
rect 207850 59520 208000 59590
rect 204000 59480 208000 59520
rect 204000 59410 204150 59480
rect 204350 59410 204650 59480
rect 204850 59410 205150 59480
rect 205350 59410 205650 59480
rect 205850 59410 206150 59480
rect 206350 59410 206650 59480
rect 206850 59410 207150 59480
rect 207350 59410 207650 59480
rect 207850 59410 208000 59480
rect 204000 59400 208000 59410
rect 204000 59380 204120 59400
rect 204380 59380 204620 59400
rect 204880 59380 205120 59400
rect 205380 59380 205620 59400
rect 205880 59380 206120 59400
rect 206380 59380 206620 59400
rect 206880 59380 207120 59400
rect 207380 59380 207620 59400
rect 207880 59380 208000 59400
rect 204000 59350 204100 59380
rect 204000 59150 204020 59350
rect 204090 59150 204100 59350
rect 204000 59120 204100 59150
rect 204400 59350 204600 59380
rect 204400 59150 204410 59350
rect 204480 59150 204520 59350
rect 204590 59150 204600 59350
rect 204400 59120 204600 59150
rect 204900 59350 205100 59380
rect 204900 59150 204910 59350
rect 204980 59150 205020 59350
rect 205090 59150 205100 59350
rect 204900 59120 205100 59150
rect 205400 59350 205600 59380
rect 205400 59150 205410 59350
rect 205480 59150 205520 59350
rect 205590 59150 205600 59350
rect 205400 59120 205600 59150
rect 205900 59350 206100 59380
rect 205900 59150 205910 59350
rect 205980 59150 206020 59350
rect 206090 59150 206100 59350
rect 205900 59120 206100 59150
rect 206400 59350 206600 59380
rect 206400 59150 206410 59350
rect 206480 59150 206520 59350
rect 206590 59150 206600 59350
rect 206400 59120 206600 59150
rect 206900 59350 207100 59380
rect 206900 59150 206910 59350
rect 206980 59150 207020 59350
rect 207090 59150 207100 59350
rect 206900 59120 207100 59150
rect 207400 59350 207600 59380
rect 207400 59150 207410 59350
rect 207480 59150 207520 59350
rect 207590 59150 207600 59350
rect 207400 59120 207600 59150
rect 207900 59350 208000 59380
rect 207900 59150 207910 59350
rect 207980 59150 208000 59350
rect 207900 59120 208000 59150
rect 204000 59100 204120 59120
rect 204380 59100 204620 59120
rect 204880 59100 205120 59120
rect 205380 59100 205620 59120
rect 205880 59100 206120 59120
rect 206380 59100 206620 59120
rect 206880 59100 207120 59120
rect 207380 59100 207620 59120
rect 207880 59100 208000 59120
rect 204000 59090 208000 59100
rect 204000 59020 204150 59090
rect 204350 59020 204650 59090
rect 204850 59020 205150 59090
rect 205350 59020 205650 59090
rect 205850 59020 206150 59090
rect 206350 59020 206650 59090
rect 206850 59020 207150 59090
rect 207350 59020 207650 59090
rect 207850 59020 208000 59090
rect 204000 58980 208000 59020
rect 204000 58910 204150 58980
rect 204350 58910 204650 58980
rect 204850 58910 205150 58980
rect 205350 58910 205650 58980
rect 205850 58910 206150 58980
rect 206350 58910 206650 58980
rect 206850 58910 207150 58980
rect 207350 58910 207650 58980
rect 207850 58910 208000 58980
rect 204000 58900 208000 58910
rect 204000 58880 204120 58900
rect 204380 58880 204620 58900
rect 204880 58880 205120 58900
rect 205380 58880 205620 58900
rect 205880 58880 206120 58900
rect 206380 58880 206620 58900
rect 206880 58880 207120 58900
rect 207380 58880 207620 58900
rect 207880 58880 208000 58900
rect 204000 58850 204100 58880
rect 204000 58650 204020 58850
rect 204090 58650 204100 58850
rect 204000 58620 204100 58650
rect 204400 58850 204600 58880
rect 204400 58650 204410 58850
rect 204480 58650 204520 58850
rect 204590 58650 204600 58850
rect 204400 58620 204600 58650
rect 204900 58850 205100 58880
rect 204900 58650 204910 58850
rect 204980 58650 205020 58850
rect 205090 58650 205100 58850
rect 204900 58620 205100 58650
rect 205400 58850 205600 58880
rect 205400 58650 205410 58850
rect 205480 58650 205520 58850
rect 205590 58650 205600 58850
rect 205400 58620 205600 58650
rect 205900 58850 206100 58880
rect 205900 58650 205910 58850
rect 205980 58650 206020 58850
rect 206090 58650 206100 58850
rect 205900 58620 206100 58650
rect 206400 58850 206600 58880
rect 206400 58650 206410 58850
rect 206480 58650 206520 58850
rect 206590 58650 206600 58850
rect 206400 58620 206600 58650
rect 206900 58850 207100 58880
rect 206900 58650 206910 58850
rect 206980 58650 207020 58850
rect 207090 58650 207100 58850
rect 206900 58620 207100 58650
rect 207400 58850 207600 58880
rect 207400 58650 207410 58850
rect 207480 58650 207520 58850
rect 207590 58650 207600 58850
rect 207400 58620 207600 58650
rect 207900 58850 208000 58880
rect 207900 58650 207910 58850
rect 207980 58650 208000 58850
rect 207900 58620 208000 58650
rect 204000 58600 204120 58620
rect 204380 58600 204620 58620
rect 204880 58600 205120 58620
rect 205380 58600 205620 58620
rect 205880 58600 206120 58620
rect 206380 58600 206620 58620
rect 206880 58600 207120 58620
rect 207380 58600 207620 58620
rect 207880 58600 208000 58620
rect 204000 58590 208000 58600
rect 204000 58520 204150 58590
rect 204350 58520 204650 58590
rect 204850 58520 205150 58590
rect 205350 58520 205650 58590
rect 205850 58520 206150 58590
rect 206350 58520 206650 58590
rect 206850 58520 207150 58590
rect 207350 58520 207650 58590
rect 207850 58520 208000 58590
rect 204000 58480 208000 58520
rect 204000 58410 204150 58480
rect 204350 58410 204650 58480
rect 204850 58410 205150 58480
rect 205350 58410 205650 58480
rect 205850 58410 206150 58480
rect 206350 58410 206650 58480
rect 206850 58410 207150 58480
rect 207350 58410 207650 58480
rect 207850 58410 208000 58480
rect 204000 58400 208000 58410
rect 204000 58380 204120 58400
rect 204380 58380 204620 58400
rect 204880 58380 205120 58400
rect 205380 58380 205620 58400
rect 205880 58380 206120 58400
rect 206380 58380 206620 58400
rect 206880 58380 207120 58400
rect 207380 58380 207620 58400
rect 207880 58380 208000 58400
rect 204000 58350 204100 58380
rect 204000 58150 204020 58350
rect 204090 58150 204100 58350
rect 204000 58120 204100 58150
rect 204400 58350 204600 58380
rect 204400 58150 204410 58350
rect 204480 58150 204520 58350
rect 204590 58150 204600 58350
rect 204400 58120 204600 58150
rect 204900 58350 205100 58380
rect 204900 58150 204910 58350
rect 204980 58150 205020 58350
rect 205090 58150 205100 58350
rect 204900 58120 205100 58150
rect 205400 58350 205600 58380
rect 205400 58150 205410 58350
rect 205480 58150 205520 58350
rect 205590 58150 205600 58350
rect 205400 58120 205600 58150
rect 205900 58350 206100 58380
rect 205900 58150 205910 58350
rect 205980 58150 206020 58350
rect 206090 58150 206100 58350
rect 205900 58120 206100 58150
rect 206400 58350 206600 58380
rect 206400 58150 206410 58350
rect 206480 58150 206520 58350
rect 206590 58150 206600 58350
rect 206400 58120 206600 58150
rect 206900 58350 207100 58380
rect 206900 58150 206910 58350
rect 206980 58150 207020 58350
rect 207090 58150 207100 58350
rect 206900 58120 207100 58150
rect 207400 58350 207600 58380
rect 207400 58150 207410 58350
rect 207480 58150 207520 58350
rect 207590 58150 207600 58350
rect 207400 58120 207600 58150
rect 207900 58350 208000 58380
rect 207900 58150 207910 58350
rect 207980 58150 208000 58350
rect 207900 58120 208000 58150
rect 204000 58100 204120 58120
rect 204380 58100 204620 58120
rect 204880 58100 205120 58120
rect 205380 58100 205620 58120
rect 205880 58100 206120 58120
rect 206380 58100 206620 58120
rect 206880 58100 207120 58120
rect 207380 58100 207620 58120
rect 207880 58100 208000 58120
rect 204000 58090 208000 58100
rect 204000 58020 204150 58090
rect 204350 58020 204650 58090
rect 204850 58020 205150 58090
rect 205350 58020 205650 58090
rect 205850 58020 206150 58090
rect 206350 58020 206650 58090
rect 206850 58020 207150 58090
rect 207350 58020 207650 58090
rect 207850 58020 208000 58090
rect 204000 57980 208000 58020
rect 204000 57910 204150 57980
rect 204350 57910 204650 57980
rect 204850 57910 205150 57980
rect 205350 57910 205650 57980
rect 205850 57910 206150 57980
rect 206350 57910 206650 57980
rect 206850 57910 207150 57980
rect 207350 57910 207650 57980
rect 207850 57910 208000 57980
rect 204000 57900 208000 57910
rect 204000 57880 204120 57900
rect 204380 57880 204620 57900
rect 204880 57880 205120 57900
rect 205380 57880 205620 57900
rect 205880 57880 206120 57900
rect 206380 57880 206620 57900
rect 206880 57880 207120 57900
rect 207380 57880 207620 57900
rect 207880 57880 208000 57900
rect 204000 57850 204100 57880
rect 204000 57650 204020 57850
rect 204090 57650 204100 57850
rect 204000 57620 204100 57650
rect 204400 57850 204600 57880
rect 204400 57650 204410 57850
rect 204480 57650 204520 57850
rect 204590 57650 204600 57850
rect 204400 57620 204600 57650
rect 204900 57850 205100 57880
rect 204900 57650 204910 57850
rect 204980 57650 205020 57850
rect 205090 57650 205100 57850
rect 204900 57620 205100 57650
rect 205400 57850 205600 57880
rect 205400 57650 205410 57850
rect 205480 57650 205520 57850
rect 205590 57650 205600 57850
rect 205400 57620 205600 57650
rect 205900 57850 206100 57880
rect 205900 57650 205910 57850
rect 205980 57650 206020 57850
rect 206090 57650 206100 57850
rect 205900 57620 206100 57650
rect 206400 57850 206600 57880
rect 206400 57650 206410 57850
rect 206480 57650 206520 57850
rect 206590 57650 206600 57850
rect 206400 57620 206600 57650
rect 206900 57850 207100 57880
rect 206900 57650 206910 57850
rect 206980 57650 207020 57850
rect 207090 57650 207100 57850
rect 206900 57620 207100 57650
rect 207400 57850 207600 57880
rect 207400 57650 207410 57850
rect 207480 57650 207520 57850
rect 207590 57650 207600 57850
rect 207400 57620 207600 57650
rect 207900 57850 208000 57880
rect 207900 57650 207910 57850
rect 207980 57650 208000 57850
rect 207900 57620 208000 57650
rect 204000 57600 204120 57620
rect 204380 57600 204620 57620
rect 204880 57600 205120 57620
rect 205380 57600 205620 57620
rect 205880 57600 206120 57620
rect 206380 57600 206620 57620
rect 206880 57600 207120 57620
rect 207380 57600 207620 57620
rect 207880 57600 208000 57620
rect 204000 57590 208000 57600
rect 204000 57520 204150 57590
rect 204350 57520 204650 57590
rect 204850 57520 205150 57590
rect 205350 57520 205650 57590
rect 205850 57520 206150 57590
rect 206350 57520 206650 57590
rect 206850 57520 207150 57590
rect 207350 57520 207650 57590
rect 207850 57520 208000 57590
rect 204000 57480 208000 57520
rect 204000 57410 204150 57480
rect 204350 57410 204650 57480
rect 204850 57410 205150 57480
rect 205350 57410 205650 57480
rect 205850 57410 206150 57480
rect 206350 57410 206650 57480
rect 206850 57410 207150 57480
rect 207350 57410 207650 57480
rect 207850 57410 208000 57480
rect 204000 57400 208000 57410
rect 204000 57380 204120 57400
rect 204380 57380 204620 57400
rect 204880 57380 205120 57400
rect 205380 57380 205620 57400
rect 205880 57380 206120 57400
rect 206380 57380 206620 57400
rect 206880 57380 207120 57400
rect 207380 57380 207620 57400
rect 207880 57380 208000 57400
rect 204000 57350 204100 57380
rect 204000 57150 204020 57350
rect 204090 57150 204100 57350
rect 204000 57120 204100 57150
rect 204400 57350 204600 57380
rect 204400 57150 204410 57350
rect 204480 57150 204520 57350
rect 204590 57150 204600 57350
rect 204400 57120 204600 57150
rect 204900 57350 205100 57380
rect 204900 57150 204910 57350
rect 204980 57150 205020 57350
rect 205090 57150 205100 57350
rect 204900 57120 205100 57150
rect 205400 57350 205600 57380
rect 205400 57150 205410 57350
rect 205480 57150 205520 57350
rect 205590 57150 205600 57350
rect 205400 57120 205600 57150
rect 205900 57350 206100 57380
rect 205900 57150 205910 57350
rect 205980 57150 206020 57350
rect 206090 57150 206100 57350
rect 205900 57120 206100 57150
rect 206400 57350 206600 57380
rect 206400 57150 206410 57350
rect 206480 57150 206520 57350
rect 206590 57150 206600 57350
rect 206400 57120 206600 57150
rect 206900 57350 207100 57380
rect 206900 57150 206910 57350
rect 206980 57150 207020 57350
rect 207090 57150 207100 57350
rect 206900 57120 207100 57150
rect 207400 57350 207600 57380
rect 207400 57150 207410 57350
rect 207480 57150 207520 57350
rect 207590 57150 207600 57350
rect 207400 57120 207600 57150
rect 207900 57350 208000 57380
rect 207900 57150 207910 57350
rect 207980 57150 208000 57350
rect 207900 57120 208000 57150
rect 204000 57100 204120 57120
rect 204380 57100 204620 57120
rect 204880 57100 205120 57120
rect 205380 57100 205620 57120
rect 205880 57100 206120 57120
rect 206380 57100 206620 57120
rect 206880 57100 207120 57120
rect 207380 57100 207620 57120
rect 207880 57100 208000 57120
rect 204000 57090 208000 57100
rect 204000 57020 204150 57090
rect 204350 57020 204650 57090
rect 204850 57020 205150 57090
rect 205350 57020 205650 57090
rect 205850 57020 206150 57090
rect 206350 57020 206650 57090
rect 206850 57020 207150 57090
rect 207350 57020 207650 57090
rect 207850 57020 208000 57090
rect 204000 56980 208000 57020
rect 204000 56910 204150 56980
rect 204350 56910 204650 56980
rect 204850 56910 205150 56980
rect 205350 56910 205650 56980
rect 205850 56910 206150 56980
rect 206350 56910 206650 56980
rect 206850 56910 207150 56980
rect 207350 56910 207650 56980
rect 207850 56910 208000 56980
rect 204000 56900 208000 56910
rect 204000 56880 204120 56900
rect 204380 56880 204620 56900
rect 204880 56880 205120 56900
rect 205380 56880 205620 56900
rect 205880 56880 206120 56900
rect 206380 56880 206620 56900
rect 206880 56880 207120 56900
rect 207380 56880 207620 56900
rect 207880 56880 208000 56900
rect 204000 56850 204100 56880
rect 204000 56650 204020 56850
rect 204090 56650 204100 56850
rect 204000 56620 204100 56650
rect 204400 56850 204600 56880
rect 204400 56650 204410 56850
rect 204480 56650 204520 56850
rect 204590 56650 204600 56850
rect 204400 56620 204600 56650
rect 204900 56850 205100 56880
rect 204900 56650 204910 56850
rect 204980 56650 205020 56850
rect 205090 56650 205100 56850
rect 204900 56620 205100 56650
rect 205400 56850 205600 56880
rect 205400 56650 205410 56850
rect 205480 56650 205520 56850
rect 205590 56650 205600 56850
rect 205400 56620 205600 56650
rect 205900 56850 206100 56880
rect 205900 56650 205910 56850
rect 205980 56650 206020 56850
rect 206090 56650 206100 56850
rect 205900 56620 206100 56650
rect 206400 56850 206600 56880
rect 206400 56650 206410 56850
rect 206480 56650 206520 56850
rect 206590 56650 206600 56850
rect 206400 56620 206600 56650
rect 206900 56850 207100 56880
rect 206900 56650 206910 56850
rect 206980 56650 207020 56850
rect 207090 56650 207100 56850
rect 206900 56620 207100 56650
rect 207400 56850 207600 56880
rect 207400 56650 207410 56850
rect 207480 56650 207520 56850
rect 207590 56650 207600 56850
rect 207400 56620 207600 56650
rect 207900 56850 208000 56880
rect 207900 56650 207910 56850
rect 207980 56650 208000 56850
rect 207900 56620 208000 56650
rect 204000 56600 204120 56620
rect 204380 56600 204620 56620
rect 204880 56600 205120 56620
rect 205380 56600 205620 56620
rect 205880 56600 206120 56620
rect 206380 56600 206620 56620
rect 206880 56600 207120 56620
rect 207380 56600 207620 56620
rect 207880 56600 208000 56620
rect 204000 56590 208000 56600
rect 204000 56520 204150 56590
rect 204350 56520 204650 56590
rect 204850 56520 205150 56590
rect 205350 56520 205650 56590
rect 205850 56520 206150 56590
rect 206350 56520 206650 56590
rect 206850 56520 207150 56590
rect 207350 56520 207650 56590
rect 207850 56520 208000 56590
rect 204000 56480 208000 56520
rect 204000 56410 204150 56480
rect 204350 56410 204650 56480
rect 204850 56410 205150 56480
rect 205350 56410 205650 56480
rect 205850 56410 206150 56480
rect 206350 56410 206650 56480
rect 206850 56410 207150 56480
rect 207350 56410 207650 56480
rect 207850 56410 208000 56480
rect 204000 56400 208000 56410
rect 204000 56380 204120 56400
rect 204380 56380 204620 56400
rect 204880 56380 205120 56400
rect 205380 56380 205620 56400
rect 205880 56380 206120 56400
rect 206380 56380 206620 56400
rect 206880 56380 207120 56400
rect 207380 56380 207620 56400
rect 207880 56380 208000 56400
rect 204000 56350 204100 56380
rect 204000 56150 204020 56350
rect 204090 56150 204100 56350
rect 204000 56120 204100 56150
rect 204400 56350 204600 56380
rect 204400 56150 204410 56350
rect 204480 56150 204520 56350
rect 204590 56150 204600 56350
rect 204400 56120 204600 56150
rect 204900 56350 205100 56380
rect 204900 56150 204910 56350
rect 204980 56150 205020 56350
rect 205090 56150 205100 56350
rect 204900 56120 205100 56150
rect 205400 56350 205600 56380
rect 205400 56150 205410 56350
rect 205480 56150 205520 56350
rect 205590 56150 205600 56350
rect 205400 56120 205600 56150
rect 205900 56350 206100 56380
rect 205900 56150 205910 56350
rect 205980 56150 206020 56350
rect 206090 56150 206100 56350
rect 205900 56120 206100 56150
rect 206400 56350 206600 56380
rect 206400 56150 206410 56350
rect 206480 56150 206520 56350
rect 206590 56150 206600 56350
rect 206400 56120 206600 56150
rect 206900 56350 207100 56380
rect 206900 56150 206910 56350
rect 206980 56150 207020 56350
rect 207090 56150 207100 56350
rect 206900 56120 207100 56150
rect 207400 56350 207600 56380
rect 207400 56150 207410 56350
rect 207480 56150 207520 56350
rect 207590 56150 207600 56350
rect 207400 56120 207600 56150
rect 207900 56350 208000 56380
rect 207900 56150 207910 56350
rect 207980 56150 208000 56350
rect 207900 56120 208000 56150
rect 204000 56100 204120 56120
rect 204380 56100 204620 56120
rect 204880 56100 205120 56120
rect 205380 56100 205620 56120
rect 205880 56100 206120 56120
rect 206380 56100 206620 56120
rect 206880 56100 207120 56120
rect 207380 56100 207620 56120
rect 207880 56100 208000 56120
rect 204000 56090 208000 56100
rect 204000 56020 204150 56090
rect 204350 56020 204650 56090
rect 204850 56020 205150 56090
rect 205350 56020 205650 56090
rect 205850 56020 206150 56090
rect 206350 56020 206650 56090
rect 206850 56020 207150 56090
rect 207350 56020 207650 56090
rect 207850 56020 208000 56090
rect 204000 55980 208000 56020
rect 204000 55910 204150 55980
rect 204350 55910 204650 55980
rect 204850 55910 205150 55980
rect 205350 55910 205650 55980
rect 205850 55910 206150 55980
rect 206350 55910 206650 55980
rect 206850 55910 207150 55980
rect 207350 55910 207650 55980
rect 207850 55910 208000 55980
rect 204000 55900 208000 55910
rect 204000 55880 204120 55900
rect 204380 55880 204620 55900
rect 204880 55880 205120 55900
rect 205380 55880 205620 55900
rect 205880 55880 206120 55900
rect 206380 55880 206620 55900
rect 206880 55880 207120 55900
rect 207380 55880 207620 55900
rect 207880 55880 208000 55900
rect 204000 55850 204100 55880
rect 204000 55650 204020 55850
rect 204090 55650 204100 55850
rect 204000 55620 204100 55650
rect 204400 55850 204600 55880
rect 204400 55650 204410 55850
rect 204480 55650 204520 55850
rect 204590 55650 204600 55850
rect 204400 55620 204600 55650
rect 204900 55850 205100 55880
rect 204900 55650 204910 55850
rect 204980 55650 205020 55850
rect 205090 55650 205100 55850
rect 204900 55620 205100 55650
rect 205400 55850 205600 55880
rect 205400 55650 205410 55850
rect 205480 55650 205520 55850
rect 205590 55650 205600 55850
rect 205400 55620 205600 55650
rect 205900 55850 206100 55880
rect 205900 55650 205910 55850
rect 205980 55650 206020 55850
rect 206090 55650 206100 55850
rect 205900 55620 206100 55650
rect 206400 55850 206600 55880
rect 206400 55650 206410 55850
rect 206480 55650 206520 55850
rect 206590 55650 206600 55850
rect 206400 55620 206600 55650
rect 206900 55850 207100 55880
rect 206900 55650 206910 55850
rect 206980 55650 207020 55850
rect 207090 55650 207100 55850
rect 206900 55620 207100 55650
rect 207400 55850 207600 55880
rect 207400 55650 207410 55850
rect 207480 55650 207520 55850
rect 207590 55650 207600 55850
rect 207400 55620 207600 55650
rect 207900 55850 208000 55880
rect 207900 55650 207910 55850
rect 207980 55650 208000 55850
rect 207900 55620 208000 55650
rect 204000 55600 204120 55620
rect 204380 55600 204620 55620
rect 204880 55600 205120 55620
rect 205380 55600 205620 55620
rect 205880 55600 206120 55620
rect 206380 55600 206620 55620
rect 206880 55600 207120 55620
rect 207380 55600 207620 55620
rect 207880 55600 208000 55620
rect 204000 55590 208000 55600
rect 204000 55520 204150 55590
rect 204350 55520 204650 55590
rect 204850 55520 205150 55590
rect 205350 55520 205650 55590
rect 205850 55520 206150 55590
rect 206350 55520 206650 55590
rect 206850 55520 207150 55590
rect 207350 55520 207650 55590
rect 207850 55520 208000 55590
rect 204000 55480 208000 55520
rect 204000 55410 204150 55480
rect 204350 55410 204650 55480
rect 204850 55410 205150 55480
rect 205350 55410 205650 55480
rect 205850 55410 206150 55480
rect 206350 55410 206650 55480
rect 206850 55410 207150 55480
rect 207350 55410 207650 55480
rect 207850 55410 208000 55480
rect 204000 55400 208000 55410
rect 204000 55380 204120 55400
rect 204380 55380 204620 55400
rect 204880 55380 205120 55400
rect 205380 55380 205620 55400
rect 205880 55380 206120 55400
rect 206380 55380 206620 55400
rect 206880 55380 207120 55400
rect 207380 55380 207620 55400
rect 207880 55380 208000 55400
rect 204000 55350 204100 55380
rect 204000 55150 204020 55350
rect 204090 55150 204100 55350
rect 204000 55120 204100 55150
rect 204400 55350 204600 55380
rect 204400 55150 204410 55350
rect 204480 55150 204520 55350
rect 204590 55150 204600 55350
rect 204400 55120 204600 55150
rect 204900 55350 205100 55380
rect 204900 55150 204910 55350
rect 204980 55150 205020 55350
rect 205090 55150 205100 55350
rect 204900 55120 205100 55150
rect 205400 55350 205600 55380
rect 205400 55150 205410 55350
rect 205480 55150 205520 55350
rect 205590 55150 205600 55350
rect 205400 55120 205600 55150
rect 205900 55350 206100 55380
rect 205900 55150 205910 55350
rect 205980 55150 206020 55350
rect 206090 55150 206100 55350
rect 205900 55120 206100 55150
rect 206400 55350 206600 55380
rect 206400 55150 206410 55350
rect 206480 55150 206520 55350
rect 206590 55150 206600 55350
rect 206400 55120 206600 55150
rect 206900 55350 207100 55380
rect 206900 55150 206910 55350
rect 206980 55150 207020 55350
rect 207090 55150 207100 55350
rect 206900 55120 207100 55150
rect 207400 55350 207600 55380
rect 207400 55150 207410 55350
rect 207480 55150 207520 55350
rect 207590 55150 207600 55350
rect 207400 55120 207600 55150
rect 207900 55350 208000 55380
rect 207900 55150 207910 55350
rect 207980 55150 208000 55350
rect 207900 55120 208000 55150
rect 204000 55100 204120 55120
rect 204380 55100 204620 55120
rect 204880 55100 205120 55120
rect 205380 55100 205620 55120
rect 205880 55100 206120 55120
rect 206380 55100 206620 55120
rect 206880 55100 207120 55120
rect 207380 55100 207620 55120
rect 207880 55100 208000 55120
rect 204000 55090 208000 55100
rect 204000 55020 204150 55090
rect 204350 55020 204650 55090
rect 204850 55020 205150 55090
rect 205350 55020 205650 55090
rect 205850 55020 206150 55090
rect 206350 55020 206650 55090
rect 206850 55020 207150 55090
rect 207350 55020 207650 55090
rect 207850 55020 208000 55090
rect 204000 54980 208000 55020
rect 204000 54910 204150 54980
rect 204350 54910 204650 54980
rect 204850 54910 205150 54980
rect 205350 54910 205650 54980
rect 205850 54910 206150 54980
rect 206350 54910 206650 54980
rect 206850 54910 207150 54980
rect 207350 54910 207650 54980
rect 207850 54910 208000 54980
rect 204000 54900 208000 54910
rect 204000 54880 204120 54900
rect 204380 54880 204620 54900
rect 204880 54880 205120 54900
rect 205380 54880 205620 54900
rect 205880 54880 206120 54900
rect 206380 54880 206620 54900
rect 206880 54880 207120 54900
rect 207380 54880 207620 54900
rect 207880 54880 208000 54900
rect 204000 54850 204100 54880
rect 204000 54650 204020 54850
rect 204090 54650 204100 54850
rect 204000 54620 204100 54650
rect 204400 54850 204600 54880
rect 204400 54650 204410 54850
rect 204480 54650 204520 54850
rect 204590 54650 204600 54850
rect 204400 54620 204600 54650
rect 204900 54850 205100 54880
rect 204900 54650 204910 54850
rect 204980 54650 205020 54850
rect 205090 54650 205100 54850
rect 204900 54620 205100 54650
rect 205400 54850 205600 54880
rect 205400 54650 205410 54850
rect 205480 54650 205520 54850
rect 205590 54650 205600 54850
rect 205400 54620 205600 54650
rect 205900 54850 206100 54880
rect 205900 54650 205910 54850
rect 205980 54650 206020 54850
rect 206090 54650 206100 54850
rect 205900 54620 206100 54650
rect 206400 54850 206600 54880
rect 206400 54650 206410 54850
rect 206480 54650 206520 54850
rect 206590 54650 206600 54850
rect 206400 54620 206600 54650
rect 206900 54850 207100 54880
rect 206900 54650 206910 54850
rect 206980 54650 207020 54850
rect 207090 54650 207100 54850
rect 206900 54620 207100 54650
rect 207400 54850 207600 54880
rect 207400 54650 207410 54850
rect 207480 54650 207520 54850
rect 207590 54650 207600 54850
rect 207400 54620 207600 54650
rect 207900 54850 208000 54880
rect 207900 54650 207910 54850
rect 207980 54650 208000 54850
rect 207900 54620 208000 54650
rect 204000 54600 204120 54620
rect 204380 54600 204620 54620
rect 204880 54600 205120 54620
rect 205380 54600 205620 54620
rect 205880 54600 206120 54620
rect 206380 54600 206620 54620
rect 206880 54600 207120 54620
rect 207380 54600 207620 54620
rect 207880 54600 208000 54620
rect 204000 54590 208000 54600
rect 204000 54520 204150 54590
rect 204350 54520 204650 54590
rect 204850 54520 205150 54590
rect 205350 54520 205650 54590
rect 205850 54520 206150 54590
rect 206350 54520 206650 54590
rect 206850 54520 207150 54590
rect 207350 54520 207650 54590
rect 207850 54520 208000 54590
rect 204000 54480 208000 54520
rect 204000 54410 204150 54480
rect 204350 54410 204650 54480
rect 204850 54410 205150 54480
rect 205350 54410 205650 54480
rect 205850 54410 206150 54480
rect 206350 54410 206650 54480
rect 206850 54410 207150 54480
rect 207350 54410 207650 54480
rect 207850 54410 208000 54480
rect 204000 54400 208000 54410
rect 204000 54380 204120 54400
rect 204380 54380 204620 54400
rect 204880 54380 205120 54400
rect 205380 54380 205620 54400
rect 205880 54380 206120 54400
rect 206380 54380 206620 54400
rect 206880 54380 207120 54400
rect 207380 54380 207620 54400
rect 207880 54380 208000 54400
rect 204000 54350 204100 54380
rect 204000 54150 204020 54350
rect 204090 54150 204100 54350
rect 204000 54120 204100 54150
rect 204400 54350 204600 54380
rect 204400 54150 204410 54350
rect 204480 54150 204520 54350
rect 204590 54150 204600 54350
rect 204400 54120 204600 54150
rect 204900 54350 205100 54380
rect 204900 54150 204910 54350
rect 204980 54150 205020 54350
rect 205090 54150 205100 54350
rect 204900 54120 205100 54150
rect 205400 54350 205600 54380
rect 205400 54150 205410 54350
rect 205480 54150 205520 54350
rect 205590 54150 205600 54350
rect 205400 54120 205600 54150
rect 205900 54350 206100 54380
rect 205900 54150 205910 54350
rect 205980 54150 206020 54350
rect 206090 54150 206100 54350
rect 205900 54120 206100 54150
rect 206400 54350 206600 54380
rect 206400 54150 206410 54350
rect 206480 54150 206520 54350
rect 206590 54150 206600 54350
rect 206400 54120 206600 54150
rect 206900 54350 207100 54380
rect 206900 54150 206910 54350
rect 206980 54150 207020 54350
rect 207090 54150 207100 54350
rect 206900 54120 207100 54150
rect 207400 54350 207600 54380
rect 207400 54150 207410 54350
rect 207480 54150 207520 54350
rect 207590 54150 207600 54350
rect 207400 54120 207600 54150
rect 207900 54350 208000 54380
rect 207900 54150 207910 54350
rect 207980 54150 208000 54350
rect 207900 54120 208000 54150
rect 204000 54100 204120 54120
rect 204380 54100 204620 54120
rect 204880 54100 205120 54120
rect 205380 54100 205620 54120
rect 205880 54100 206120 54120
rect 206380 54100 206620 54120
rect 206880 54100 207120 54120
rect 207380 54100 207620 54120
rect 207880 54100 208000 54120
rect 204000 54090 208000 54100
rect 204000 54020 204150 54090
rect 204350 54020 204650 54090
rect 204850 54020 205150 54090
rect 205350 54020 205650 54090
rect 205850 54020 206150 54090
rect 206350 54020 206650 54090
rect 206850 54020 207150 54090
rect 207350 54020 207650 54090
rect 207850 54020 208000 54090
rect 204000 53980 208000 54020
rect 204000 53910 204150 53980
rect 204350 53910 204650 53980
rect 204850 53910 205150 53980
rect 205350 53910 205650 53980
rect 205850 53910 206150 53980
rect 206350 53910 206650 53980
rect 206850 53910 207150 53980
rect 207350 53910 207650 53980
rect 207850 53910 208000 53980
rect 204000 53900 208000 53910
rect 204000 53880 204120 53900
rect 204380 53880 204620 53900
rect 204880 53880 205120 53900
rect 205380 53880 205620 53900
rect 205880 53880 206120 53900
rect 206380 53880 206620 53900
rect 206880 53880 207120 53900
rect 207380 53880 207620 53900
rect 207880 53880 208000 53900
rect 204000 53850 204100 53880
rect 204000 53650 204020 53850
rect 204090 53650 204100 53850
rect 204000 53620 204100 53650
rect 204400 53850 204600 53880
rect 204400 53650 204410 53850
rect 204480 53650 204520 53850
rect 204590 53650 204600 53850
rect 204400 53620 204600 53650
rect 204900 53850 205100 53880
rect 204900 53650 204910 53850
rect 204980 53650 205020 53850
rect 205090 53650 205100 53850
rect 204900 53620 205100 53650
rect 205400 53850 205600 53880
rect 205400 53650 205410 53850
rect 205480 53650 205520 53850
rect 205590 53650 205600 53850
rect 205400 53620 205600 53650
rect 205900 53850 206100 53880
rect 205900 53650 205910 53850
rect 205980 53650 206020 53850
rect 206090 53650 206100 53850
rect 205900 53620 206100 53650
rect 206400 53850 206600 53880
rect 206400 53650 206410 53850
rect 206480 53650 206520 53850
rect 206590 53650 206600 53850
rect 206400 53620 206600 53650
rect 206900 53850 207100 53880
rect 206900 53650 206910 53850
rect 206980 53650 207020 53850
rect 207090 53650 207100 53850
rect 206900 53620 207100 53650
rect 207400 53850 207600 53880
rect 207400 53650 207410 53850
rect 207480 53650 207520 53850
rect 207590 53650 207600 53850
rect 207400 53620 207600 53650
rect 207900 53850 208000 53880
rect 207900 53650 207910 53850
rect 207980 53650 208000 53850
rect 207900 53620 208000 53650
rect 204000 53600 204120 53620
rect 204380 53600 204620 53620
rect 204880 53600 205120 53620
rect 205380 53600 205620 53620
rect 205880 53600 206120 53620
rect 206380 53600 206620 53620
rect 206880 53600 207120 53620
rect 207380 53600 207620 53620
rect 207880 53600 208000 53620
rect 204000 53590 208000 53600
rect 204000 53520 204150 53590
rect 204350 53520 204650 53590
rect 204850 53520 205150 53590
rect 205350 53520 205650 53590
rect 205850 53520 206150 53590
rect 206350 53520 206650 53590
rect 206850 53520 207150 53590
rect 207350 53520 207650 53590
rect 207850 53520 208000 53590
rect 204000 53480 208000 53520
rect 204000 53410 204150 53480
rect 204350 53410 204650 53480
rect 204850 53410 205150 53480
rect 205350 53410 205650 53480
rect 205850 53410 206150 53480
rect 206350 53410 206650 53480
rect 206850 53410 207150 53480
rect 207350 53410 207650 53480
rect 207850 53410 208000 53480
rect 204000 53400 208000 53410
rect 204000 53380 204120 53400
rect 204380 53380 204620 53400
rect 204880 53380 205120 53400
rect 205380 53380 205620 53400
rect 205880 53380 206120 53400
rect 206380 53380 206620 53400
rect 206880 53380 207120 53400
rect 207380 53380 207620 53400
rect 207880 53380 208000 53400
rect 204000 53350 204100 53380
rect 204000 53150 204020 53350
rect 204090 53150 204100 53350
rect 204000 53120 204100 53150
rect 204400 53350 204600 53380
rect 204400 53150 204410 53350
rect 204480 53150 204520 53350
rect 204590 53150 204600 53350
rect 204400 53120 204600 53150
rect 204900 53350 205100 53380
rect 204900 53150 204910 53350
rect 204980 53150 205020 53350
rect 205090 53150 205100 53350
rect 204900 53120 205100 53150
rect 205400 53350 205600 53380
rect 205400 53150 205410 53350
rect 205480 53150 205520 53350
rect 205590 53150 205600 53350
rect 205400 53120 205600 53150
rect 205900 53350 206100 53380
rect 205900 53150 205910 53350
rect 205980 53150 206020 53350
rect 206090 53150 206100 53350
rect 205900 53120 206100 53150
rect 206400 53350 206600 53380
rect 206400 53150 206410 53350
rect 206480 53150 206520 53350
rect 206590 53150 206600 53350
rect 206400 53120 206600 53150
rect 206900 53350 207100 53380
rect 206900 53150 206910 53350
rect 206980 53150 207020 53350
rect 207090 53150 207100 53350
rect 206900 53120 207100 53150
rect 207400 53350 207600 53380
rect 207400 53150 207410 53350
rect 207480 53150 207520 53350
rect 207590 53150 207600 53350
rect 207400 53120 207600 53150
rect 207900 53350 208000 53380
rect 207900 53150 207910 53350
rect 207980 53150 208000 53350
rect 207900 53120 208000 53150
rect 204000 53100 204120 53120
rect 204380 53100 204620 53120
rect 204880 53100 205120 53120
rect 205380 53100 205620 53120
rect 205880 53100 206120 53120
rect 206380 53100 206620 53120
rect 206880 53100 207120 53120
rect 207380 53100 207620 53120
rect 207880 53100 208000 53120
rect 204000 53090 208000 53100
rect 204000 53020 204150 53090
rect 204350 53020 204650 53090
rect 204850 53020 205150 53090
rect 205350 53020 205650 53090
rect 205850 53020 206150 53090
rect 206350 53020 206650 53090
rect 206850 53020 207150 53090
rect 207350 53020 207650 53090
rect 207850 53020 208000 53090
rect 204000 52980 208000 53020
rect 204000 52910 204150 52980
rect 204350 52910 204650 52980
rect 204850 52910 205150 52980
rect 205350 52910 205650 52980
rect 205850 52910 206150 52980
rect 206350 52910 206650 52980
rect 206850 52910 207150 52980
rect 207350 52910 207650 52980
rect 207850 52910 208000 52980
rect 204000 52900 208000 52910
rect 204000 52880 204120 52900
rect 204380 52880 204620 52900
rect 204880 52880 205120 52900
rect 205380 52880 205620 52900
rect 205880 52880 206120 52900
rect 206380 52880 206620 52900
rect 206880 52880 207120 52900
rect 207380 52880 207620 52900
rect 207880 52880 208000 52900
rect 204000 52850 204100 52880
rect 204000 52650 204020 52850
rect 204090 52650 204100 52850
rect 204000 52620 204100 52650
rect 204400 52850 204600 52880
rect 204400 52650 204410 52850
rect 204480 52650 204520 52850
rect 204590 52650 204600 52850
rect 204400 52620 204600 52650
rect 204900 52850 205100 52880
rect 204900 52650 204910 52850
rect 204980 52650 205020 52850
rect 205090 52650 205100 52850
rect 204900 52620 205100 52650
rect 205400 52850 205600 52880
rect 205400 52650 205410 52850
rect 205480 52650 205520 52850
rect 205590 52650 205600 52850
rect 205400 52620 205600 52650
rect 205900 52850 206100 52880
rect 205900 52650 205910 52850
rect 205980 52650 206020 52850
rect 206090 52650 206100 52850
rect 205900 52620 206100 52650
rect 206400 52850 206600 52880
rect 206400 52650 206410 52850
rect 206480 52650 206520 52850
rect 206590 52650 206600 52850
rect 206400 52620 206600 52650
rect 206900 52850 207100 52880
rect 206900 52650 206910 52850
rect 206980 52650 207020 52850
rect 207090 52650 207100 52850
rect 206900 52620 207100 52650
rect 207400 52850 207600 52880
rect 207400 52650 207410 52850
rect 207480 52650 207520 52850
rect 207590 52650 207600 52850
rect 207400 52620 207600 52650
rect 207900 52850 208000 52880
rect 207900 52650 207910 52850
rect 207980 52650 208000 52850
rect 207900 52620 208000 52650
rect 204000 52600 204120 52620
rect 204380 52600 204620 52620
rect 204880 52600 205120 52620
rect 205380 52600 205620 52620
rect 205880 52600 206120 52620
rect 206380 52600 206620 52620
rect 206880 52600 207120 52620
rect 207380 52600 207620 52620
rect 207880 52600 208000 52620
rect 204000 52590 208000 52600
rect 204000 52520 204150 52590
rect 204350 52520 204650 52590
rect 204850 52520 205150 52590
rect 205350 52520 205650 52590
rect 205850 52520 206150 52590
rect 206350 52520 206650 52590
rect 206850 52520 207150 52590
rect 207350 52520 207650 52590
rect 207850 52520 208000 52590
rect 204000 52480 208000 52520
rect 204000 52410 204150 52480
rect 204350 52410 204650 52480
rect 204850 52410 205150 52480
rect 205350 52410 205650 52480
rect 205850 52410 206150 52480
rect 206350 52410 206650 52480
rect 206850 52410 207150 52480
rect 207350 52410 207650 52480
rect 207850 52410 208000 52480
rect 204000 52400 208000 52410
rect 204000 52380 204120 52400
rect 204380 52380 204620 52400
rect 204880 52380 205120 52400
rect 205380 52380 205620 52400
rect 205880 52380 206120 52400
rect 206380 52380 206620 52400
rect 206880 52380 207120 52400
rect 207380 52380 207620 52400
rect 207880 52380 208000 52400
rect 204000 52350 204100 52380
rect 204000 52150 204020 52350
rect 204090 52150 204100 52350
rect 204000 52120 204100 52150
rect 204400 52350 204600 52380
rect 204400 52150 204410 52350
rect 204480 52150 204520 52350
rect 204590 52150 204600 52350
rect 204400 52120 204600 52150
rect 204900 52350 205100 52380
rect 204900 52150 204910 52350
rect 204980 52150 205020 52350
rect 205090 52150 205100 52350
rect 204900 52120 205100 52150
rect 205400 52350 205600 52380
rect 205400 52150 205410 52350
rect 205480 52150 205520 52350
rect 205590 52150 205600 52350
rect 205400 52120 205600 52150
rect 205900 52350 206100 52380
rect 205900 52150 205910 52350
rect 205980 52150 206020 52350
rect 206090 52150 206100 52350
rect 205900 52120 206100 52150
rect 206400 52350 206600 52380
rect 206400 52150 206410 52350
rect 206480 52150 206520 52350
rect 206590 52150 206600 52350
rect 206400 52120 206600 52150
rect 206900 52350 207100 52380
rect 206900 52150 206910 52350
rect 206980 52150 207020 52350
rect 207090 52150 207100 52350
rect 206900 52120 207100 52150
rect 207400 52350 207600 52380
rect 207400 52150 207410 52350
rect 207480 52150 207520 52350
rect 207590 52150 207600 52350
rect 207400 52120 207600 52150
rect 207900 52350 208000 52380
rect 207900 52150 207910 52350
rect 207980 52150 208000 52350
rect 207900 52120 208000 52150
rect 204000 52100 204120 52120
rect 204380 52100 204620 52120
rect 204880 52100 205120 52120
rect 205380 52100 205620 52120
rect 205880 52100 206120 52120
rect 206380 52100 206620 52120
rect 206880 52100 207120 52120
rect 207380 52100 207620 52120
rect 207880 52100 208000 52120
rect 204000 52090 208000 52100
rect 204000 52020 204150 52090
rect 204350 52020 204650 52090
rect 204850 52020 205150 52090
rect 205350 52020 205650 52090
rect 205850 52020 206150 52090
rect 206350 52020 206650 52090
rect 206850 52020 207150 52090
rect 207350 52020 207650 52090
rect 207850 52020 208000 52090
rect 204000 51980 208000 52020
rect 204000 51910 204150 51980
rect 204350 51910 204650 51980
rect 204850 51910 205150 51980
rect 205350 51910 205650 51980
rect 205850 51910 206150 51980
rect 206350 51910 206650 51980
rect 206850 51910 207150 51980
rect 207350 51910 207650 51980
rect 207850 51910 208000 51980
rect 204000 51900 208000 51910
rect 204000 51880 204120 51900
rect 204380 51880 204620 51900
rect 204880 51880 205120 51900
rect 205380 51880 205620 51900
rect 205880 51880 206120 51900
rect 206380 51880 206620 51900
rect 206880 51880 207120 51900
rect 207380 51880 207620 51900
rect 207880 51880 208000 51900
rect 204000 51850 204100 51880
rect 204000 51650 204020 51850
rect 204090 51650 204100 51850
rect 204000 51620 204100 51650
rect 204400 51850 204600 51880
rect 204400 51650 204410 51850
rect 204480 51650 204520 51850
rect 204590 51650 204600 51850
rect 204400 51620 204600 51650
rect 204900 51850 205100 51880
rect 204900 51650 204910 51850
rect 204980 51650 205020 51850
rect 205090 51650 205100 51850
rect 204900 51620 205100 51650
rect 205400 51850 205600 51880
rect 205400 51650 205410 51850
rect 205480 51650 205520 51850
rect 205590 51650 205600 51850
rect 205400 51620 205600 51650
rect 205900 51850 206100 51880
rect 205900 51650 205910 51850
rect 205980 51650 206020 51850
rect 206090 51650 206100 51850
rect 205900 51620 206100 51650
rect 206400 51850 206600 51880
rect 206400 51650 206410 51850
rect 206480 51650 206520 51850
rect 206590 51650 206600 51850
rect 206400 51620 206600 51650
rect 206900 51850 207100 51880
rect 206900 51650 206910 51850
rect 206980 51650 207020 51850
rect 207090 51650 207100 51850
rect 206900 51620 207100 51650
rect 207400 51850 207600 51880
rect 207400 51650 207410 51850
rect 207480 51650 207520 51850
rect 207590 51650 207600 51850
rect 207400 51620 207600 51650
rect 207900 51850 208000 51880
rect 207900 51650 207910 51850
rect 207980 51650 208000 51850
rect 207900 51620 208000 51650
rect 204000 51600 204120 51620
rect 204380 51600 204620 51620
rect 204880 51600 205120 51620
rect 205380 51600 205620 51620
rect 205880 51600 206120 51620
rect 206380 51600 206620 51620
rect 206880 51600 207120 51620
rect 207380 51600 207620 51620
rect 207880 51600 208000 51620
rect 204000 51590 208000 51600
rect 204000 51520 204150 51590
rect 204350 51520 204650 51590
rect 204850 51520 205150 51590
rect 205350 51520 205650 51590
rect 205850 51520 206150 51590
rect 206350 51520 206650 51590
rect 206850 51520 207150 51590
rect 207350 51520 207650 51590
rect 207850 51520 208000 51590
rect 204000 51480 208000 51520
rect 204000 51410 204150 51480
rect 204350 51410 204650 51480
rect 204850 51410 205150 51480
rect 205350 51410 205650 51480
rect 205850 51410 206150 51480
rect 206350 51410 206650 51480
rect 206850 51410 207150 51480
rect 207350 51410 207650 51480
rect 207850 51410 208000 51480
rect 204000 51400 208000 51410
rect 204000 51380 204120 51400
rect 204380 51380 204620 51400
rect 204880 51380 205120 51400
rect 205380 51380 205620 51400
rect 205880 51380 206120 51400
rect 206380 51380 206620 51400
rect 206880 51380 207120 51400
rect 207380 51380 207620 51400
rect 207880 51380 208000 51400
rect 204000 51350 204100 51380
rect 204000 51150 204020 51350
rect 204090 51150 204100 51350
rect 204000 51120 204100 51150
rect 204400 51350 204600 51380
rect 204400 51150 204410 51350
rect 204480 51150 204520 51350
rect 204590 51150 204600 51350
rect 204400 51120 204600 51150
rect 204900 51350 205100 51380
rect 204900 51150 204910 51350
rect 204980 51150 205020 51350
rect 205090 51150 205100 51350
rect 204900 51120 205100 51150
rect 205400 51350 205600 51380
rect 205400 51150 205410 51350
rect 205480 51150 205520 51350
rect 205590 51150 205600 51350
rect 205400 51120 205600 51150
rect 205900 51350 206100 51380
rect 205900 51150 205910 51350
rect 205980 51150 206020 51350
rect 206090 51150 206100 51350
rect 205900 51120 206100 51150
rect 206400 51350 206600 51380
rect 206400 51150 206410 51350
rect 206480 51150 206520 51350
rect 206590 51150 206600 51350
rect 206400 51120 206600 51150
rect 206900 51350 207100 51380
rect 206900 51150 206910 51350
rect 206980 51150 207020 51350
rect 207090 51150 207100 51350
rect 206900 51120 207100 51150
rect 207400 51350 207600 51380
rect 207400 51150 207410 51350
rect 207480 51150 207520 51350
rect 207590 51150 207600 51350
rect 207400 51120 207600 51150
rect 207900 51350 208000 51380
rect 207900 51150 207910 51350
rect 207980 51150 208000 51350
rect 207900 51120 208000 51150
rect 204000 51100 204120 51120
rect 204380 51100 204620 51120
rect 204880 51100 205120 51120
rect 205380 51100 205620 51120
rect 205880 51100 206120 51120
rect 206380 51100 206620 51120
rect 206880 51100 207120 51120
rect 207380 51100 207620 51120
rect 207880 51100 208000 51120
rect 204000 51090 208000 51100
rect 204000 51020 204150 51090
rect 204350 51020 204650 51090
rect 204850 51020 205150 51090
rect 205350 51020 205650 51090
rect 205850 51020 206150 51090
rect 206350 51020 206650 51090
rect 206850 51020 207150 51090
rect 207350 51020 207650 51090
rect 207850 51020 208000 51090
rect 204000 50980 208000 51020
rect 204000 50910 204150 50980
rect 204350 50910 204650 50980
rect 204850 50910 205150 50980
rect 205350 50910 205650 50980
rect 205850 50910 206150 50980
rect 206350 50910 206650 50980
rect 206850 50910 207150 50980
rect 207350 50910 207650 50980
rect 207850 50910 208000 50980
rect 204000 50900 208000 50910
rect 204000 50880 204120 50900
rect 204380 50880 204620 50900
rect 204880 50880 205120 50900
rect 205380 50880 205620 50900
rect 205880 50880 206120 50900
rect 206380 50880 206620 50900
rect 206880 50880 207120 50900
rect 207380 50880 207620 50900
rect 207880 50880 208000 50900
rect 204000 50850 204100 50880
rect 204000 50650 204020 50850
rect 204090 50650 204100 50850
rect 204000 50620 204100 50650
rect 204400 50850 204600 50880
rect 204400 50650 204410 50850
rect 204480 50650 204520 50850
rect 204590 50650 204600 50850
rect 204400 50620 204600 50650
rect 204900 50850 205100 50880
rect 204900 50650 204910 50850
rect 204980 50650 205020 50850
rect 205090 50650 205100 50850
rect 204900 50620 205100 50650
rect 205400 50850 205600 50880
rect 205400 50650 205410 50850
rect 205480 50650 205520 50850
rect 205590 50650 205600 50850
rect 205400 50620 205600 50650
rect 205900 50850 206100 50880
rect 205900 50650 205910 50850
rect 205980 50650 206020 50850
rect 206090 50650 206100 50850
rect 205900 50620 206100 50650
rect 206400 50850 206600 50880
rect 206400 50650 206410 50850
rect 206480 50650 206520 50850
rect 206590 50650 206600 50850
rect 206400 50620 206600 50650
rect 206900 50850 207100 50880
rect 206900 50650 206910 50850
rect 206980 50650 207020 50850
rect 207090 50650 207100 50850
rect 206900 50620 207100 50650
rect 207400 50850 207600 50880
rect 207400 50650 207410 50850
rect 207480 50650 207520 50850
rect 207590 50650 207600 50850
rect 207400 50620 207600 50650
rect 207900 50850 208000 50880
rect 207900 50650 207910 50850
rect 207980 50650 208000 50850
rect 207900 50620 208000 50650
rect 204000 50600 204120 50620
rect 204380 50600 204620 50620
rect 204880 50600 205120 50620
rect 205380 50600 205620 50620
rect 205880 50600 206120 50620
rect 206380 50600 206620 50620
rect 206880 50600 207120 50620
rect 207380 50600 207620 50620
rect 207880 50600 208000 50620
rect 204000 50590 208000 50600
rect 204000 50520 204150 50590
rect 204350 50520 204650 50590
rect 204850 50520 205150 50590
rect 205350 50520 205650 50590
rect 205850 50520 206150 50590
rect 206350 50520 206650 50590
rect 206850 50520 207150 50590
rect 207350 50520 207650 50590
rect 207850 50520 208000 50590
rect 204000 50480 208000 50520
rect 204000 50410 204150 50480
rect 204350 50410 204650 50480
rect 204850 50410 205150 50480
rect 205350 50410 205650 50480
rect 205850 50410 206150 50480
rect 206350 50410 206650 50480
rect 206850 50410 207150 50480
rect 207350 50410 207650 50480
rect 207850 50410 208000 50480
rect 204000 50400 208000 50410
rect 204000 50380 204120 50400
rect 204380 50380 204620 50400
rect 204880 50380 205120 50400
rect 205380 50380 205620 50400
rect 205880 50380 206120 50400
rect 206380 50380 206620 50400
rect 206880 50380 207120 50400
rect 207380 50380 207620 50400
rect 207880 50380 208000 50400
rect 204000 50350 204100 50380
rect 204000 50150 204020 50350
rect 204090 50150 204100 50350
rect 204000 50120 204100 50150
rect 204400 50350 204600 50380
rect 204400 50150 204410 50350
rect 204480 50150 204520 50350
rect 204590 50150 204600 50350
rect 204400 50120 204600 50150
rect 204900 50350 205100 50380
rect 204900 50150 204910 50350
rect 204980 50150 205020 50350
rect 205090 50150 205100 50350
rect 204900 50120 205100 50150
rect 205400 50350 205600 50380
rect 205400 50150 205410 50350
rect 205480 50150 205520 50350
rect 205590 50150 205600 50350
rect 205400 50120 205600 50150
rect 205900 50350 206100 50380
rect 205900 50150 205910 50350
rect 205980 50150 206020 50350
rect 206090 50150 206100 50350
rect 205900 50120 206100 50150
rect 206400 50350 206600 50380
rect 206400 50150 206410 50350
rect 206480 50150 206520 50350
rect 206590 50150 206600 50350
rect 206400 50120 206600 50150
rect 206900 50350 207100 50380
rect 206900 50150 206910 50350
rect 206980 50150 207020 50350
rect 207090 50150 207100 50350
rect 206900 50120 207100 50150
rect 207400 50350 207600 50380
rect 207400 50150 207410 50350
rect 207480 50150 207520 50350
rect 207590 50150 207600 50350
rect 207400 50120 207600 50150
rect 207900 50350 208000 50380
rect 207900 50150 207910 50350
rect 207980 50150 208000 50350
rect 207900 50120 208000 50150
rect 204000 50100 204120 50120
rect 204380 50100 204620 50120
rect 204880 50100 205120 50120
rect 205380 50100 205620 50120
rect 205880 50100 206120 50120
rect 206380 50100 206620 50120
rect 206880 50100 207120 50120
rect 207380 50100 207620 50120
rect 207880 50100 208000 50120
rect 204000 50090 208000 50100
rect 204000 50020 204150 50090
rect 204350 50020 204650 50090
rect 204850 50020 205150 50090
rect 205350 50020 205650 50090
rect 205850 50020 206150 50090
rect 206350 50020 206650 50090
rect 206850 50020 207150 50090
rect 207350 50020 207650 50090
rect 207850 50020 208000 50090
rect 204000 49980 208000 50020
rect 204000 49910 204150 49980
rect 204350 49910 204650 49980
rect 204850 49910 205150 49980
rect 205350 49910 205650 49980
rect 205850 49910 206150 49980
rect 206350 49910 206650 49980
rect 206850 49910 207150 49980
rect 207350 49910 207650 49980
rect 207850 49910 208000 49980
rect 204000 49900 208000 49910
rect 204000 49880 204120 49900
rect 204380 49880 204620 49900
rect 204880 49880 205120 49900
rect 205380 49880 205620 49900
rect 205880 49880 206120 49900
rect 206380 49880 206620 49900
rect 206880 49880 207120 49900
rect 207380 49880 207620 49900
rect 207880 49880 208000 49900
rect 204000 49850 204100 49880
rect 204000 49650 204020 49850
rect 204090 49650 204100 49850
rect 204000 49620 204100 49650
rect 204400 49850 204600 49880
rect 204400 49650 204410 49850
rect 204480 49650 204520 49850
rect 204590 49650 204600 49850
rect 204400 49620 204600 49650
rect 204900 49850 205100 49880
rect 204900 49650 204910 49850
rect 204980 49650 205020 49850
rect 205090 49650 205100 49850
rect 204900 49620 205100 49650
rect 205400 49850 205600 49880
rect 205400 49650 205410 49850
rect 205480 49650 205520 49850
rect 205590 49650 205600 49850
rect 205400 49620 205600 49650
rect 205900 49850 206100 49880
rect 205900 49650 205910 49850
rect 205980 49650 206020 49850
rect 206090 49650 206100 49850
rect 205900 49620 206100 49650
rect 206400 49850 206600 49880
rect 206400 49650 206410 49850
rect 206480 49650 206520 49850
rect 206590 49650 206600 49850
rect 206400 49620 206600 49650
rect 206900 49850 207100 49880
rect 206900 49650 206910 49850
rect 206980 49650 207020 49850
rect 207090 49650 207100 49850
rect 206900 49620 207100 49650
rect 207400 49850 207600 49880
rect 207400 49650 207410 49850
rect 207480 49650 207520 49850
rect 207590 49650 207600 49850
rect 207400 49620 207600 49650
rect 207900 49850 208000 49880
rect 207900 49650 207910 49850
rect 207980 49650 208000 49850
rect 207900 49620 208000 49650
rect 204000 49600 204120 49620
rect 204380 49600 204620 49620
rect 204880 49600 205120 49620
rect 205380 49600 205620 49620
rect 205880 49600 206120 49620
rect 206380 49600 206620 49620
rect 206880 49600 207120 49620
rect 207380 49600 207620 49620
rect 207880 49600 208000 49620
rect 204000 49590 208000 49600
rect 204000 49520 204150 49590
rect 204350 49520 204650 49590
rect 204850 49520 205150 49590
rect 205350 49520 205650 49590
rect 205850 49520 206150 49590
rect 206350 49520 206650 49590
rect 206850 49520 207150 49590
rect 207350 49520 207650 49590
rect 207850 49520 208000 49590
rect 204000 49480 208000 49520
rect 204000 49410 204150 49480
rect 204350 49410 204650 49480
rect 204850 49410 205150 49480
rect 205350 49410 205650 49480
rect 205850 49410 206150 49480
rect 206350 49410 206650 49480
rect 206850 49410 207150 49480
rect 207350 49410 207650 49480
rect 207850 49410 208000 49480
rect 204000 49400 208000 49410
rect 204000 49380 204120 49400
rect 204380 49380 204620 49400
rect 204880 49380 205120 49400
rect 205380 49380 205620 49400
rect 205880 49380 206120 49400
rect 206380 49380 206620 49400
rect 206880 49380 207120 49400
rect 207380 49380 207620 49400
rect 207880 49380 208000 49400
rect 204000 49350 204100 49380
rect 204000 49150 204020 49350
rect 204090 49150 204100 49350
rect 204000 49120 204100 49150
rect 204400 49350 204600 49380
rect 204400 49150 204410 49350
rect 204480 49150 204520 49350
rect 204590 49150 204600 49350
rect 204400 49120 204600 49150
rect 204900 49350 205100 49380
rect 204900 49150 204910 49350
rect 204980 49150 205020 49350
rect 205090 49150 205100 49350
rect 204900 49120 205100 49150
rect 205400 49350 205600 49380
rect 205400 49150 205410 49350
rect 205480 49150 205520 49350
rect 205590 49150 205600 49350
rect 205400 49120 205600 49150
rect 205900 49350 206100 49380
rect 205900 49150 205910 49350
rect 205980 49150 206020 49350
rect 206090 49150 206100 49350
rect 205900 49120 206100 49150
rect 206400 49350 206600 49380
rect 206400 49150 206410 49350
rect 206480 49150 206520 49350
rect 206590 49150 206600 49350
rect 206400 49120 206600 49150
rect 206900 49350 207100 49380
rect 206900 49150 206910 49350
rect 206980 49150 207020 49350
rect 207090 49150 207100 49350
rect 206900 49120 207100 49150
rect 207400 49350 207600 49380
rect 207400 49150 207410 49350
rect 207480 49150 207520 49350
rect 207590 49150 207600 49350
rect 207400 49120 207600 49150
rect 207900 49350 208000 49380
rect 207900 49150 207910 49350
rect 207980 49150 208000 49350
rect 207900 49120 208000 49150
rect 204000 49100 204120 49120
rect 204380 49100 204620 49120
rect 204880 49100 205120 49120
rect 205380 49100 205620 49120
rect 205880 49100 206120 49120
rect 206380 49100 206620 49120
rect 206880 49100 207120 49120
rect 207380 49100 207620 49120
rect 207880 49100 208000 49120
rect 204000 49090 208000 49100
rect 204000 49020 204150 49090
rect 204350 49020 204650 49090
rect 204850 49020 205150 49090
rect 205350 49020 205650 49090
rect 205850 49020 206150 49090
rect 206350 49020 206650 49090
rect 206850 49020 207150 49090
rect 207350 49020 207650 49090
rect 207850 49020 208000 49090
rect 204000 48980 208000 49020
rect 204000 48910 204150 48980
rect 204350 48910 204650 48980
rect 204850 48910 205150 48980
rect 205350 48910 205650 48980
rect 205850 48910 206150 48980
rect 206350 48910 206650 48980
rect 206850 48910 207150 48980
rect 207350 48910 207650 48980
rect 207850 48910 208000 48980
rect 204000 48900 208000 48910
rect 204000 48880 204120 48900
rect 204380 48880 204620 48900
rect 204880 48880 205120 48900
rect 205380 48880 205620 48900
rect 205880 48880 206120 48900
rect 206380 48880 206620 48900
rect 206880 48880 207120 48900
rect 207380 48880 207620 48900
rect 207880 48880 208000 48900
rect 204000 48850 204100 48880
rect 204000 48650 204020 48850
rect 204090 48650 204100 48850
rect 204000 48620 204100 48650
rect 204400 48850 204600 48880
rect 204400 48650 204410 48850
rect 204480 48650 204520 48850
rect 204590 48650 204600 48850
rect 204400 48620 204600 48650
rect 204900 48850 205100 48880
rect 204900 48650 204910 48850
rect 204980 48650 205020 48850
rect 205090 48650 205100 48850
rect 204900 48620 205100 48650
rect 205400 48850 205600 48880
rect 205400 48650 205410 48850
rect 205480 48650 205520 48850
rect 205590 48650 205600 48850
rect 205400 48620 205600 48650
rect 205900 48850 206100 48880
rect 205900 48650 205910 48850
rect 205980 48650 206020 48850
rect 206090 48650 206100 48850
rect 205900 48620 206100 48650
rect 206400 48850 206600 48880
rect 206400 48650 206410 48850
rect 206480 48650 206520 48850
rect 206590 48650 206600 48850
rect 206400 48620 206600 48650
rect 206900 48850 207100 48880
rect 206900 48650 206910 48850
rect 206980 48650 207020 48850
rect 207090 48650 207100 48850
rect 206900 48620 207100 48650
rect 207400 48850 207600 48880
rect 207400 48650 207410 48850
rect 207480 48650 207520 48850
rect 207590 48650 207600 48850
rect 207400 48620 207600 48650
rect 207900 48850 208000 48880
rect 207900 48650 207910 48850
rect 207980 48650 208000 48850
rect 207900 48620 208000 48650
rect 204000 48600 204120 48620
rect 204380 48600 204620 48620
rect 204880 48600 205120 48620
rect 205380 48600 205620 48620
rect 205880 48600 206120 48620
rect 206380 48600 206620 48620
rect 206880 48600 207120 48620
rect 207380 48600 207620 48620
rect 207880 48600 208000 48620
rect 204000 48590 208000 48600
rect 204000 48520 204150 48590
rect 204350 48520 204650 48590
rect 204850 48520 205150 48590
rect 205350 48520 205650 48590
rect 205850 48520 206150 48590
rect 206350 48520 206650 48590
rect 206850 48520 207150 48590
rect 207350 48520 207650 48590
rect 207850 48520 208000 48590
rect 204000 48480 208000 48520
rect 204000 48410 204150 48480
rect 204350 48410 204650 48480
rect 204850 48410 205150 48480
rect 205350 48410 205650 48480
rect 205850 48410 206150 48480
rect 206350 48410 206650 48480
rect 206850 48410 207150 48480
rect 207350 48410 207650 48480
rect 207850 48410 208000 48480
rect 204000 48400 208000 48410
rect 204000 48380 204120 48400
rect 204380 48380 204620 48400
rect 204880 48380 205120 48400
rect 205380 48380 205620 48400
rect 205880 48380 206120 48400
rect 206380 48380 206620 48400
rect 206880 48380 207120 48400
rect 207380 48380 207620 48400
rect 207880 48380 208000 48400
rect 204000 48350 204100 48380
rect 204000 48150 204020 48350
rect 204090 48150 204100 48350
rect 204000 48120 204100 48150
rect 204400 48350 204600 48380
rect 204400 48150 204410 48350
rect 204480 48150 204520 48350
rect 204590 48150 204600 48350
rect 204400 48120 204600 48150
rect 204900 48350 205100 48380
rect 204900 48150 204910 48350
rect 204980 48150 205020 48350
rect 205090 48150 205100 48350
rect 204900 48120 205100 48150
rect 205400 48350 205600 48380
rect 205400 48150 205410 48350
rect 205480 48150 205520 48350
rect 205590 48150 205600 48350
rect 205400 48120 205600 48150
rect 205900 48350 206100 48380
rect 205900 48150 205910 48350
rect 205980 48150 206020 48350
rect 206090 48150 206100 48350
rect 205900 48120 206100 48150
rect 206400 48350 206600 48380
rect 206400 48150 206410 48350
rect 206480 48150 206520 48350
rect 206590 48150 206600 48350
rect 206400 48120 206600 48150
rect 206900 48350 207100 48380
rect 206900 48150 206910 48350
rect 206980 48150 207020 48350
rect 207090 48150 207100 48350
rect 206900 48120 207100 48150
rect 207400 48350 207600 48380
rect 207400 48150 207410 48350
rect 207480 48150 207520 48350
rect 207590 48150 207600 48350
rect 207400 48120 207600 48150
rect 207900 48350 208000 48380
rect 207900 48150 207910 48350
rect 207980 48150 208000 48350
rect 207900 48120 208000 48150
rect 204000 48100 204120 48120
rect 204380 48100 204620 48120
rect 204880 48100 205120 48120
rect 205380 48100 205620 48120
rect 205880 48100 206120 48120
rect 206380 48100 206620 48120
rect 206880 48100 207120 48120
rect 207380 48100 207620 48120
rect 207880 48100 208000 48120
rect 204000 48090 208000 48100
rect 204000 48020 204150 48090
rect 204350 48020 204650 48090
rect 204850 48020 205150 48090
rect 205350 48020 205650 48090
rect 205850 48020 206150 48090
rect 206350 48020 206650 48090
rect 206850 48020 207150 48090
rect 207350 48020 207650 48090
rect 207850 48020 208000 48090
rect 204000 47980 208000 48020
rect 204000 47910 204150 47980
rect 204350 47910 204650 47980
rect 204850 47910 205150 47980
rect 205350 47910 205650 47980
rect 205850 47910 206150 47980
rect 206350 47910 206650 47980
rect 206850 47910 207150 47980
rect 207350 47910 207650 47980
rect 207850 47910 208000 47980
rect 204000 47900 208000 47910
rect 204000 47880 204120 47900
rect 204380 47880 204620 47900
rect 204880 47880 205120 47900
rect 205380 47880 205620 47900
rect 205880 47880 206120 47900
rect 206380 47880 206620 47900
rect 206880 47880 207120 47900
rect 207380 47880 207620 47900
rect 207880 47880 208000 47900
rect 204000 47850 204100 47880
rect 204000 47650 204020 47850
rect 204090 47650 204100 47850
rect 204000 47620 204100 47650
rect 204400 47850 204600 47880
rect 204400 47650 204410 47850
rect 204480 47650 204520 47850
rect 204590 47650 204600 47850
rect 204400 47620 204600 47650
rect 204900 47850 205100 47880
rect 204900 47650 204910 47850
rect 204980 47650 205020 47850
rect 205090 47650 205100 47850
rect 204900 47620 205100 47650
rect 205400 47850 205600 47880
rect 205400 47650 205410 47850
rect 205480 47650 205520 47850
rect 205590 47650 205600 47850
rect 205400 47620 205600 47650
rect 205900 47850 206100 47880
rect 205900 47650 205910 47850
rect 205980 47650 206020 47850
rect 206090 47650 206100 47850
rect 205900 47620 206100 47650
rect 206400 47850 206600 47880
rect 206400 47650 206410 47850
rect 206480 47650 206520 47850
rect 206590 47650 206600 47850
rect 206400 47620 206600 47650
rect 206900 47850 207100 47880
rect 206900 47650 206910 47850
rect 206980 47650 207020 47850
rect 207090 47650 207100 47850
rect 206900 47620 207100 47650
rect 207400 47850 207600 47880
rect 207400 47650 207410 47850
rect 207480 47650 207520 47850
rect 207590 47650 207600 47850
rect 207400 47620 207600 47650
rect 207900 47850 208000 47880
rect 207900 47650 207910 47850
rect 207980 47650 208000 47850
rect 207900 47620 208000 47650
rect 204000 47600 204120 47620
rect 204380 47600 204620 47620
rect 204880 47600 205120 47620
rect 205380 47600 205620 47620
rect 205880 47600 206120 47620
rect 206380 47600 206620 47620
rect 206880 47600 207120 47620
rect 207380 47600 207620 47620
rect 207880 47600 208000 47620
rect 204000 47590 208000 47600
rect 204000 47520 204150 47590
rect 204350 47520 204650 47590
rect 204850 47520 205150 47590
rect 205350 47520 205650 47590
rect 205850 47520 206150 47590
rect 206350 47520 206650 47590
rect 206850 47520 207150 47590
rect 207350 47520 207650 47590
rect 207850 47520 208000 47590
rect 204000 47480 208000 47520
rect 204000 47410 204150 47480
rect 204350 47410 204650 47480
rect 204850 47410 205150 47480
rect 205350 47410 205650 47480
rect 205850 47410 206150 47480
rect 206350 47410 206650 47480
rect 206850 47410 207150 47480
rect 207350 47410 207650 47480
rect 207850 47410 208000 47480
rect 204000 47400 208000 47410
rect 204000 47380 204120 47400
rect 204380 47380 204620 47400
rect 204880 47380 205120 47400
rect 205380 47380 205620 47400
rect 205880 47380 206120 47400
rect 206380 47380 206620 47400
rect 206880 47380 207120 47400
rect 207380 47380 207620 47400
rect 207880 47380 208000 47400
rect 204000 47350 204100 47380
rect 204000 47150 204020 47350
rect 204090 47150 204100 47350
rect 204000 47120 204100 47150
rect 204400 47350 204600 47380
rect 204400 47150 204410 47350
rect 204480 47150 204520 47350
rect 204590 47150 204600 47350
rect 204400 47120 204600 47150
rect 204900 47350 205100 47380
rect 204900 47150 204910 47350
rect 204980 47150 205020 47350
rect 205090 47150 205100 47350
rect 204900 47120 205100 47150
rect 205400 47350 205600 47380
rect 205400 47150 205410 47350
rect 205480 47150 205520 47350
rect 205590 47150 205600 47350
rect 205400 47120 205600 47150
rect 205900 47350 206100 47380
rect 205900 47150 205910 47350
rect 205980 47150 206020 47350
rect 206090 47150 206100 47350
rect 205900 47120 206100 47150
rect 206400 47350 206600 47380
rect 206400 47150 206410 47350
rect 206480 47150 206520 47350
rect 206590 47150 206600 47350
rect 206400 47120 206600 47150
rect 206900 47350 207100 47380
rect 206900 47150 206910 47350
rect 206980 47150 207020 47350
rect 207090 47150 207100 47350
rect 206900 47120 207100 47150
rect 207400 47350 207600 47380
rect 207400 47150 207410 47350
rect 207480 47150 207520 47350
rect 207590 47150 207600 47350
rect 207400 47120 207600 47150
rect 207900 47350 208000 47380
rect 207900 47150 207910 47350
rect 207980 47150 208000 47350
rect 207900 47120 208000 47150
rect 204000 47100 204120 47120
rect 204380 47100 204620 47120
rect 204880 47100 205120 47120
rect 205380 47100 205620 47120
rect 205880 47100 206120 47120
rect 206380 47100 206620 47120
rect 206880 47100 207120 47120
rect 207380 47100 207620 47120
rect 207880 47100 208000 47120
rect 204000 47090 208000 47100
rect 204000 47020 204150 47090
rect 204350 47020 204650 47090
rect 204850 47020 205150 47090
rect 205350 47020 205650 47090
rect 205850 47020 206150 47090
rect 206350 47020 206650 47090
rect 206850 47020 207150 47090
rect 207350 47020 207650 47090
rect 207850 47020 208000 47090
rect 204000 46980 208000 47020
rect 204000 46910 204150 46980
rect 204350 46910 204650 46980
rect 204850 46910 205150 46980
rect 205350 46910 205650 46980
rect 205850 46910 206150 46980
rect 206350 46910 206650 46980
rect 206850 46910 207150 46980
rect 207350 46910 207650 46980
rect 207850 46910 208000 46980
rect 204000 46900 208000 46910
rect 204000 46880 204120 46900
rect 204380 46880 204620 46900
rect 204880 46880 205120 46900
rect 205380 46880 205620 46900
rect 205880 46880 206120 46900
rect 206380 46880 206620 46900
rect 206880 46880 207120 46900
rect 207380 46880 207620 46900
rect 207880 46880 208000 46900
rect 204000 46850 204100 46880
rect 204000 46650 204020 46850
rect 204090 46650 204100 46850
rect 204000 46620 204100 46650
rect 204400 46850 204600 46880
rect 204400 46650 204410 46850
rect 204480 46650 204520 46850
rect 204590 46650 204600 46850
rect 204400 46620 204600 46650
rect 204900 46850 205100 46880
rect 204900 46650 204910 46850
rect 204980 46650 205020 46850
rect 205090 46650 205100 46850
rect 204900 46620 205100 46650
rect 205400 46850 205600 46880
rect 205400 46650 205410 46850
rect 205480 46650 205520 46850
rect 205590 46650 205600 46850
rect 205400 46620 205600 46650
rect 205900 46850 206100 46880
rect 205900 46650 205910 46850
rect 205980 46650 206020 46850
rect 206090 46650 206100 46850
rect 205900 46620 206100 46650
rect 206400 46850 206600 46880
rect 206400 46650 206410 46850
rect 206480 46650 206520 46850
rect 206590 46650 206600 46850
rect 206400 46620 206600 46650
rect 206900 46850 207100 46880
rect 206900 46650 206910 46850
rect 206980 46650 207020 46850
rect 207090 46650 207100 46850
rect 206900 46620 207100 46650
rect 207400 46850 207600 46880
rect 207400 46650 207410 46850
rect 207480 46650 207520 46850
rect 207590 46650 207600 46850
rect 207400 46620 207600 46650
rect 207900 46850 208000 46880
rect 207900 46650 207910 46850
rect 207980 46650 208000 46850
rect 207900 46620 208000 46650
rect 204000 46600 204120 46620
rect 204380 46600 204620 46620
rect 204880 46600 205120 46620
rect 205380 46600 205620 46620
rect 205880 46600 206120 46620
rect 206380 46600 206620 46620
rect 206880 46600 207120 46620
rect 207380 46600 207620 46620
rect 207880 46600 208000 46620
rect 204000 46590 208000 46600
rect 204000 46520 204150 46590
rect 204350 46520 204650 46590
rect 204850 46520 205150 46590
rect 205350 46520 205650 46590
rect 205850 46520 206150 46590
rect 206350 46520 206650 46590
rect 206850 46520 207150 46590
rect 207350 46520 207650 46590
rect 207850 46520 208000 46590
rect 204000 46480 208000 46520
rect 204000 46410 204150 46480
rect 204350 46410 204650 46480
rect 204850 46410 205150 46480
rect 205350 46410 205650 46480
rect 205850 46410 206150 46480
rect 206350 46410 206650 46480
rect 206850 46410 207150 46480
rect 207350 46410 207650 46480
rect 207850 46410 208000 46480
rect 204000 46400 208000 46410
rect 204000 46380 204120 46400
rect 204380 46380 204620 46400
rect 204880 46380 205120 46400
rect 205380 46380 205620 46400
rect 205880 46380 206120 46400
rect 206380 46380 206620 46400
rect 206880 46380 207120 46400
rect 207380 46380 207620 46400
rect 207880 46380 208000 46400
rect 204000 46350 204100 46380
rect 204000 46150 204020 46350
rect 204090 46150 204100 46350
rect 204000 46120 204100 46150
rect 204400 46350 204600 46380
rect 204400 46150 204410 46350
rect 204480 46150 204520 46350
rect 204590 46150 204600 46350
rect 204400 46120 204600 46150
rect 204900 46350 205100 46380
rect 204900 46150 204910 46350
rect 204980 46150 205020 46350
rect 205090 46150 205100 46350
rect 204900 46120 205100 46150
rect 205400 46350 205600 46380
rect 205400 46150 205410 46350
rect 205480 46150 205520 46350
rect 205590 46150 205600 46350
rect 205400 46120 205600 46150
rect 205900 46350 206100 46380
rect 205900 46150 205910 46350
rect 205980 46150 206020 46350
rect 206090 46150 206100 46350
rect 205900 46120 206100 46150
rect 206400 46350 206600 46380
rect 206400 46150 206410 46350
rect 206480 46150 206520 46350
rect 206590 46150 206600 46350
rect 206400 46120 206600 46150
rect 206900 46350 207100 46380
rect 206900 46150 206910 46350
rect 206980 46150 207020 46350
rect 207090 46150 207100 46350
rect 206900 46120 207100 46150
rect 207400 46350 207600 46380
rect 207400 46150 207410 46350
rect 207480 46150 207520 46350
rect 207590 46150 207600 46350
rect 207400 46120 207600 46150
rect 207900 46350 208000 46380
rect 207900 46150 207910 46350
rect 207980 46150 208000 46350
rect 207900 46120 208000 46150
rect 204000 46100 204120 46120
rect 204380 46100 204620 46120
rect 204880 46100 205120 46120
rect 205380 46100 205620 46120
rect 205880 46100 206120 46120
rect 206380 46100 206620 46120
rect 206880 46100 207120 46120
rect 207380 46100 207620 46120
rect 207880 46100 208000 46120
rect 204000 46090 208000 46100
rect 204000 46020 204150 46090
rect 204350 46020 204650 46090
rect 204850 46020 205150 46090
rect 205350 46020 205650 46090
rect 205850 46020 206150 46090
rect 206350 46020 206650 46090
rect 206850 46020 207150 46090
rect 207350 46020 207650 46090
rect 207850 46020 208000 46090
rect 204000 45980 208000 46020
rect 204000 45910 204150 45980
rect 204350 45910 204650 45980
rect 204850 45910 205150 45980
rect 205350 45910 205650 45980
rect 205850 45910 206150 45980
rect 206350 45910 206650 45980
rect 206850 45910 207150 45980
rect 207350 45910 207650 45980
rect 207850 45910 208000 45980
rect 204000 45900 208000 45910
rect 204000 45880 204120 45900
rect 204380 45880 204620 45900
rect 204880 45880 205120 45900
rect 205380 45880 205620 45900
rect 205880 45880 206120 45900
rect 206380 45880 206620 45900
rect 206880 45880 207120 45900
rect 207380 45880 207620 45900
rect 207880 45880 208000 45900
rect 204000 45850 204100 45880
rect 204000 45650 204020 45850
rect 204090 45650 204100 45850
rect 204000 45620 204100 45650
rect 204400 45850 204600 45880
rect 204400 45650 204410 45850
rect 204480 45650 204520 45850
rect 204590 45650 204600 45850
rect 204400 45620 204600 45650
rect 204900 45850 205100 45880
rect 204900 45650 204910 45850
rect 204980 45650 205020 45850
rect 205090 45650 205100 45850
rect 204900 45620 205100 45650
rect 205400 45850 205600 45880
rect 205400 45650 205410 45850
rect 205480 45650 205520 45850
rect 205590 45650 205600 45850
rect 205400 45620 205600 45650
rect 205900 45850 206100 45880
rect 205900 45650 205910 45850
rect 205980 45650 206020 45850
rect 206090 45650 206100 45850
rect 205900 45620 206100 45650
rect 206400 45850 206600 45880
rect 206400 45650 206410 45850
rect 206480 45650 206520 45850
rect 206590 45650 206600 45850
rect 206400 45620 206600 45650
rect 206900 45850 207100 45880
rect 206900 45650 206910 45850
rect 206980 45650 207020 45850
rect 207090 45650 207100 45850
rect 206900 45620 207100 45650
rect 207400 45850 207600 45880
rect 207400 45650 207410 45850
rect 207480 45650 207520 45850
rect 207590 45650 207600 45850
rect 207400 45620 207600 45650
rect 207900 45850 208000 45880
rect 207900 45650 207910 45850
rect 207980 45650 208000 45850
rect 207900 45620 208000 45650
rect 204000 45600 204120 45620
rect 204380 45600 204620 45620
rect 204880 45600 205120 45620
rect 205380 45600 205620 45620
rect 205880 45600 206120 45620
rect 206380 45600 206620 45620
rect 206880 45600 207120 45620
rect 207380 45600 207620 45620
rect 207880 45600 208000 45620
rect 204000 45590 208000 45600
rect 204000 45520 204150 45590
rect 204350 45520 204650 45590
rect 204850 45520 205150 45590
rect 205350 45520 205650 45590
rect 205850 45520 206150 45590
rect 206350 45520 206650 45590
rect 206850 45520 207150 45590
rect 207350 45520 207650 45590
rect 207850 45520 208000 45590
rect 204000 45480 208000 45520
rect 204000 45410 204150 45480
rect 204350 45410 204650 45480
rect 204850 45410 205150 45480
rect 205350 45410 205650 45480
rect 205850 45410 206150 45480
rect 206350 45410 206650 45480
rect 206850 45410 207150 45480
rect 207350 45410 207650 45480
rect 207850 45410 208000 45480
rect 204000 45400 208000 45410
rect 204000 45380 204120 45400
rect 204380 45380 204620 45400
rect 204880 45380 205120 45400
rect 205380 45380 205620 45400
rect 205880 45380 206120 45400
rect 206380 45380 206620 45400
rect 206880 45380 207120 45400
rect 207380 45380 207620 45400
rect 207880 45380 208000 45400
rect 204000 45350 204100 45380
rect 204000 45150 204020 45350
rect 204090 45150 204100 45350
rect 204000 45120 204100 45150
rect 204400 45350 204600 45380
rect 204400 45150 204410 45350
rect 204480 45150 204520 45350
rect 204590 45150 204600 45350
rect 204400 45120 204600 45150
rect 204900 45350 205100 45380
rect 204900 45150 204910 45350
rect 204980 45150 205020 45350
rect 205090 45150 205100 45350
rect 204900 45120 205100 45150
rect 205400 45350 205600 45380
rect 205400 45150 205410 45350
rect 205480 45150 205520 45350
rect 205590 45150 205600 45350
rect 205400 45120 205600 45150
rect 205900 45350 206100 45380
rect 205900 45150 205910 45350
rect 205980 45150 206020 45350
rect 206090 45150 206100 45350
rect 205900 45120 206100 45150
rect 206400 45350 206600 45380
rect 206400 45150 206410 45350
rect 206480 45150 206520 45350
rect 206590 45150 206600 45350
rect 206400 45120 206600 45150
rect 206900 45350 207100 45380
rect 206900 45150 206910 45350
rect 206980 45150 207020 45350
rect 207090 45150 207100 45350
rect 206900 45120 207100 45150
rect 207400 45350 207600 45380
rect 207400 45150 207410 45350
rect 207480 45150 207520 45350
rect 207590 45150 207600 45350
rect 207400 45120 207600 45150
rect 207900 45350 208000 45380
rect 207900 45150 207910 45350
rect 207980 45150 208000 45350
rect 207900 45120 208000 45150
rect 204000 45100 204120 45120
rect 204380 45100 204620 45120
rect 204880 45100 205120 45120
rect 205380 45100 205620 45120
rect 205880 45100 206120 45120
rect 206380 45100 206620 45120
rect 206880 45100 207120 45120
rect 207380 45100 207620 45120
rect 207880 45100 208000 45120
rect 204000 45090 208000 45100
rect 204000 45020 204150 45090
rect 204350 45020 204650 45090
rect 204850 45020 205150 45090
rect 205350 45020 205650 45090
rect 205850 45020 206150 45090
rect 206350 45020 206650 45090
rect 206850 45020 207150 45090
rect 207350 45020 207650 45090
rect 207850 45020 208000 45090
rect 204000 44980 208000 45020
rect 204000 44910 204150 44980
rect 204350 44910 204650 44980
rect 204850 44910 205150 44980
rect 205350 44910 205650 44980
rect 205850 44910 206150 44980
rect 206350 44910 206650 44980
rect 206850 44910 207150 44980
rect 207350 44910 207650 44980
rect 207850 44910 208000 44980
rect 204000 44900 208000 44910
rect 204000 44880 204120 44900
rect 204380 44880 204620 44900
rect 204880 44880 205120 44900
rect 205380 44880 205620 44900
rect 205880 44880 206120 44900
rect 206380 44880 206620 44900
rect 206880 44880 207120 44900
rect 207380 44880 207620 44900
rect 207880 44880 208000 44900
rect 204000 44850 204100 44880
rect 204000 44650 204020 44850
rect 204090 44650 204100 44850
rect 204000 44620 204100 44650
rect 204400 44850 204600 44880
rect 204400 44650 204410 44850
rect 204480 44650 204520 44850
rect 204590 44650 204600 44850
rect 204400 44620 204600 44650
rect 204900 44850 205100 44880
rect 204900 44650 204910 44850
rect 204980 44650 205020 44850
rect 205090 44650 205100 44850
rect 204900 44620 205100 44650
rect 205400 44850 205600 44880
rect 205400 44650 205410 44850
rect 205480 44650 205520 44850
rect 205590 44650 205600 44850
rect 205400 44620 205600 44650
rect 205900 44850 206100 44880
rect 205900 44650 205910 44850
rect 205980 44650 206020 44850
rect 206090 44650 206100 44850
rect 205900 44620 206100 44650
rect 206400 44850 206600 44880
rect 206400 44650 206410 44850
rect 206480 44650 206520 44850
rect 206590 44650 206600 44850
rect 206400 44620 206600 44650
rect 206900 44850 207100 44880
rect 206900 44650 206910 44850
rect 206980 44650 207020 44850
rect 207090 44650 207100 44850
rect 206900 44620 207100 44650
rect 207400 44850 207600 44880
rect 207400 44650 207410 44850
rect 207480 44650 207520 44850
rect 207590 44650 207600 44850
rect 207400 44620 207600 44650
rect 207900 44850 208000 44880
rect 207900 44650 207910 44850
rect 207980 44650 208000 44850
rect 207900 44620 208000 44650
rect 204000 44600 204120 44620
rect 204380 44600 204620 44620
rect 204880 44600 205120 44620
rect 205380 44600 205620 44620
rect 205880 44600 206120 44620
rect 206380 44600 206620 44620
rect 206880 44600 207120 44620
rect 207380 44600 207620 44620
rect 207880 44600 208000 44620
rect 204000 44590 208000 44600
rect 204000 44520 204150 44590
rect 204350 44520 204650 44590
rect 204850 44520 205150 44590
rect 205350 44520 205650 44590
rect 205850 44520 206150 44590
rect 206350 44520 206650 44590
rect 206850 44520 207150 44590
rect 207350 44520 207650 44590
rect 207850 44520 208000 44590
rect 204000 44480 208000 44520
rect 204000 44410 204150 44480
rect 204350 44410 204650 44480
rect 204850 44410 205150 44480
rect 205350 44410 205650 44480
rect 205850 44410 206150 44480
rect 206350 44410 206650 44480
rect 206850 44410 207150 44480
rect 207350 44410 207650 44480
rect 207850 44410 208000 44480
rect 204000 44400 208000 44410
rect 204000 44380 204120 44400
rect 204380 44380 204620 44400
rect 204880 44380 205120 44400
rect 205380 44380 205620 44400
rect 205880 44380 206120 44400
rect 206380 44380 206620 44400
rect 206880 44380 207120 44400
rect 207380 44380 207620 44400
rect 207880 44380 208000 44400
rect 204000 44350 204100 44380
rect 204000 44150 204020 44350
rect 204090 44150 204100 44350
rect 204000 44120 204100 44150
rect 204400 44350 204600 44380
rect 204400 44150 204410 44350
rect 204480 44150 204520 44350
rect 204590 44150 204600 44350
rect 204400 44120 204600 44150
rect 204900 44350 205100 44380
rect 204900 44150 204910 44350
rect 204980 44150 205020 44350
rect 205090 44150 205100 44350
rect 204900 44120 205100 44150
rect 205400 44350 205600 44380
rect 205400 44150 205410 44350
rect 205480 44150 205520 44350
rect 205590 44150 205600 44350
rect 205400 44120 205600 44150
rect 205900 44350 206100 44380
rect 205900 44150 205910 44350
rect 205980 44150 206020 44350
rect 206090 44150 206100 44350
rect 205900 44120 206100 44150
rect 206400 44350 206600 44380
rect 206400 44150 206410 44350
rect 206480 44150 206520 44350
rect 206590 44150 206600 44350
rect 206400 44120 206600 44150
rect 206900 44350 207100 44380
rect 206900 44150 206910 44350
rect 206980 44150 207020 44350
rect 207090 44150 207100 44350
rect 206900 44120 207100 44150
rect 207400 44350 207600 44380
rect 207400 44150 207410 44350
rect 207480 44150 207520 44350
rect 207590 44150 207600 44350
rect 207400 44120 207600 44150
rect 207900 44350 208000 44380
rect 207900 44150 207910 44350
rect 207980 44150 208000 44350
rect 207900 44120 208000 44150
rect 204000 44100 204120 44120
rect 204380 44100 204620 44120
rect 204880 44100 205120 44120
rect 205380 44100 205620 44120
rect 205880 44100 206120 44120
rect 206380 44100 206620 44120
rect 206880 44100 207120 44120
rect 207380 44100 207620 44120
rect 207880 44100 208000 44120
rect 204000 44090 208000 44100
rect 204000 44020 204150 44090
rect 204350 44020 204650 44090
rect 204850 44020 205150 44090
rect 205350 44020 205650 44090
rect 205850 44020 206150 44090
rect 206350 44020 206650 44090
rect 206850 44020 207150 44090
rect 207350 44020 207650 44090
rect 207850 44020 208000 44090
rect 204000 43980 208000 44020
rect 204000 43910 204150 43980
rect 204350 43910 204650 43980
rect 204850 43910 205150 43980
rect 205350 43910 205650 43980
rect 205850 43910 206150 43980
rect 206350 43910 206650 43980
rect 206850 43910 207150 43980
rect 207350 43910 207650 43980
rect 207850 43910 208000 43980
rect 204000 43900 208000 43910
rect 204000 43880 204120 43900
rect 204380 43880 204620 43900
rect 204880 43880 205120 43900
rect 205380 43880 205620 43900
rect 205880 43880 206120 43900
rect 206380 43880 206620 43900
rect 206880 43880 207120 43900
rect 207380 43880 207620 43900
rect 207880 43880 208000 43900
rect 204000 43850 204100 43880
rect 204000 43650 204020 43850
rect 204090 43650 204100 43850
rect 204000 43620 204100 43650
rect 204400 43850 204600 43880
rect 204400 43650 204410 43850
rect 204480 43650 204520 43850
rect 204590 43650 204600 43850
rect 204400 43620 204600 43650
rect 204900 43850 205100 43880
rect 204900 43650 204910 43850
rect 204980 43650 205020 43850
rect 205090 43650 205100 43850
rect 204900 43620 205100 43650
rect 205400 43850 205600 43880
rect 205400 43650 205410 43850
rect 205480 43650 205520 43850
rect 205590 43650 205600 43850
rect 205400 43620 205600 43650
rect 205900 43850 206100 43880
rect 205900 43650 205910 43850
rect 205980 43650 206020 43850
rect 206090 43650 206100 43850
rect 205900 43620 206100 43650
rect 206400 43850 206600 43880
rect 206400 43650 206410 43850
rect 206480 43650 206520 43850
rect 206590 43650 206600 43850
rect 206400 43620 206600 43650
rect 206900 43850 207100 43880
rect 206900 43650 206910 43850
rect 206980 43650 207020 43850
rect 207090 43650 207100 43850
rect 206900 43620 207100 43650
rect 207400 43850 207600 43880
rect 207400 43650 207410 43850
rect 207480 43650 207520 43850
rect 207590 43650 207600 43850
rect 207400 43620 207600 43650
rect 207900 43850 208000 43880
rect 207900 43650 207910 43850
rect 207980 43650 208000 43850
rect 207900 43620 208000 43650
rect 204000 43600 204120 43620
rect 204380 43600 204620 43620
rect 204880 43600 205120 43620
rect 205380 43600 205620 43620
rect 205880 43600 206120 43620
rect 206380 43600 206620 43620
rect 206880 43600 207120 43620
rect 207380 43600 207620 43620
rect 207880 43600 208000 43620
rect 204000 43590 208000 43600
rect 204000 43520 204150 43590
rect 204350 43520 204650 43590
rect 204850 43520 205150 43590
rect 205350 43520 205650 43590
rect 205850 43520 206150 43590
rect 206350 43520 206650 43590
rect 206850 43520 207150 43590
rect 207350 43520 207650 43590
rect 207850 43520 208000 43590
rect 204000 43480 208000 43520
rect 204000 43410 204150 43480
rect 204350 43410 204650 43480
rect 204850 43410 205150 43480
rect 205350 43410 205650 43480
rect 205850 43410 206150 43480
rect 206350 43410 206650 43480
rect 206850 43410 207150 43480
rect 207350 43410 207650 43480
rect 207850 43410 208000 43480
rect 204000 43400 208000 43410
rect 204000 43380 204120 43400
rect 204380 43380 204620 43400
rect 204880 43380 205120 43400
rect 205380 43380 205620 43400
rect 205880 43380 206120 43400
rect 206380 43380 206620 43400
rect 206880 43380 207120 43400
rect 207380 43380 207620 43400
rect 207880 43380 208000 43400
rect 204000 43350 204100 43380
rect 204000 43150 204020 43350
rect 204090 43150 204100 43350
rect 204000 43120 204100 43150
rect 204400 43350 204600 43380
rect 204400 43150 204410 43350
rect 204480 43150 204520 43350
rect 204590 43150 204600 43350
rect 204400 43120 204600 43150
rect 204900 43350 205100 43380
rect 204900 43150 204910 43350
rect 204980 43150 205020 43350
rect 205090 43150 205100 43350
rect 204900 43120 205100 43150
rect 205400 43350 205600 43380
rect 205400 43150 205410 43350
rect 205480 43150 205520 43350
rect 205590 43150 205600 43350
rect 205400 43120 205600 43150
rect 205900 43350 206100 43380
rect 205900 43150 205910 43350
rect 205980 43150 206020 43350
rect 206090 43150 206100 43350
rect 205900 43120 206100 43150
rect 206400 43350 206600 43380
rect 206400 43150 206410 43350
rect 206480 43150 206520 43350
rect 206590 43150 206600 43350
rect 206400 43120 206600 43150
rect 206900 43350 207100 43380
rect 206900 43150 206910 43350
rect 206980 43150 207020 43350
rect 207090 43150 207100 43350
rect 206900 43120 207100 43150
rect 207400 43350 207600 43380
rect 207400 43150 207410 43350
rect 207480 43150 207520 43350
rect 207590 43150 207600 43350
rect 207400 43120 207600 43150
rect 207900 43350 208000 43380
rect 207900 43150 207910 43350
rect 207980 43150 208000 43350
rect 207900 43120 208000 43150
rect 204000 43100 204120 43120
rect 204380 43100 204620 43120
rect 204880 43100 205120 43120
rect 205380 43100 205620 43120
rect 205880 43100 206120 43120
rect 206380 43100 206620 43120
rect 206880 43100 207120 43120
rect 207380 43100 207620 43120
rect 207880 43100 208000 43120
rect 204000 43090 208000 43100
rect 204000 43020 204150 43090
rect 204350 43020 204650 43090
rect 204850 43020 205150 43090
rect 205350 43020 205650 43090
rect 205850 43020 206150 43090
rect 206350 43020 206650 43090
rect 206850 43020 207150 43090
rect 207350 43020 207650 43090
rect 207850 43020 208000 43090
rect 204000 42980 208000 43020
rect 204000 42910 204150 42980
rect 204350 42910 204650 42980
rect 204850 42910 205150 42980
rect 205350 42910 205650 42980
rect 205850 42910 206150 42980
rect 206350 42910 206650 42980
rect 206850 42910 207150 42980
rect 207350 42910 207650 42980
rect 207850 42910 208000 42980
rect 204000 42900 208000 42910
rect 204000 42880 204120 42900
rect 204380 42880 204620 42900
rect 204880 42880 205120 42900
rect 205380 42880 205620 42900
rect 205880 42880 206120 42900
rect 206380 42880 206620 42900
rect 206880 42880 207120 42900
rect 207380 42880 207620 42900
rect 207880 42880 208000 42900
rect 204000 42850 204100 42880
rect 204000 42650 204020 42850
rect 204090 42650 204100 42850
rect 204000 42620 204100 42650
rect 204400 42850 204600 42880
rect 204400 42650 204410 42850
rect 204480 42650 204520 42850
rect 204590 42650 204600 42850
rect 204400 42620 204600 42650
rect 204900 42850 205100 42880
rect 204900 42650 204910 42850
rect 204980 42650 205020 42850
rect 205090 42650 205100 42850
rect 204900 42620 205100 42650
rect 205400 42850 205600 42880
rect 205400 42650 205410 42850
rect 205480 42650 205520 42850
rect 205590 42650 205600 42850
rect 205400 42620 205600 42650
rect 205900 42850 206100 42880
rect 205900 42650 205910 42850
rect 205980 42650 206020 42850
rect 206090 42650 206100 42850
rect 205900 42620 206100 42650
rect 206400 42850 206600 42880
rect 206400 42650 206410 42850
rect 206480 42650 206520 42850
rect 206590 42650 206600 42850
rect 206400 42620 206600 42650
rect 206900 42850 207100 42880
rect 206900 42650 206910 42850
rect 206980 42650 207020 42850
rect 207090 42650 207100 42850
rect 206900 42620 207100 42650
rect 207400 42850 207600 42880
rect 207400 42650 207410 42850
rect 207480 42650 207520 42850
rect 207590 42650 207600 42850
rect 207400 42620 207600 42650
rect 207900 42850 208000 42880
rect 207900 42650 207910 42850
rect 207980 42650 208000 42850
rect 207900 42620 208000 42650
rect 204000 42600 204120 42620
rect 204380 42600 204620 42620
rect 204880 42600 205120 42620
rect 205380 42600 205620 42620
rect 205880 42600 206120 42620
rect 206380 42600 206620 42620
rect 206880 42600 207120 42620
rect 207380 42600 207620 42620
rect 207880 42600 208000 42620
rect 204000 42590 208000 42600
rect 204000 42520 204150 42590
rect 204350 42520 204650 42590
rect 204850 42520 205150 42590
rect 205350 42520 205650 42590
rect 205850 42520 206150 42590
rect 206350 42520 206650 42590
rect 206850 42520 207150 42590
rect 207350 42520 207650 42590
rect 207850 42520 208000 42590
rect 204000 42480 208000 42520
rect 204000 42410 204150 42480
rect 204350 42410 204650 42480
rect 204850 42410 205150 42480
rect 205350 42410 205650 42480
rect 205850 42410 206150 42480
rect 206350 42410 206650 42480
rect 206850 42410 207150 42480
rect 207350 42410 207650 42480
rect 207850 42410 208000 42480
rect 204000 42400 208000 42410
rect 204000 42380 204120 42400
rect 204380 42380 204620 42400
rect 204880 42380 205120 42400
rect 205380 42380 205620 42400
rect 205880 42380 206120 42400
rect 206380 42380 206620 42400
rect 206880 42380 207120 42400
rect 207380 42380 207620 42400
rect 207880 42380 208000 42400
rect 204000 42350 204100 42380
rect 204000 42150 204020 42350
rect 204090 42150 204100 42350
rect 204000 42120 204100 42150
rect 204400 42350 204600 42380
rect 204400 42150 204410 42350
rect 204480 42150 204520 42350
rect 204590 42150 204600 42350
rect 204400 42120 204600 42150
rect 204900 42350 205100 42380
rect 204900 42150 204910 42350
rect 204980 42150 205020 42350
rect 205090 42150 205100 42350
rect 204900 42120 205100 42150
rect 205400 42350 205600 42380
rect 205400 42150 205410 42350
rect 205480 42150 205520 42350
rect 205590 42150 205600 42350
rect 205400 42120 205600 42150
rect 205900 42350 206100 42380
rect 205900 42150 205910 42350
rect 205980 42150 206020 42350
rect 206090 42150 206100 42350
rect 205900 42120 206100 42150
rect 206400 42350 206600 42380
rect 206400 42150 206410 42350
rect 206480 42150 206520 42350
rect 206590 42150 206600 42350
rect 206400 42120 206600 42150
rect 206900 42350 207100 42380
rect 206900 42150 206910 42350
rect 206980 42150 207020 42350
rect 207090 42150 207100 42350
rect 206900 42120 207100 42150
rect 207400 42350 207600 42380
rect 207400 42150 207410 42350
rect 207480 42150 207520 42350
rect 207590 42150 207600 42350
rect 207400 42120 207600 42150
rect 207900 42350 208000 42380
rect 207900 42150 207910 42350
rect 207980 42150 208000 42350
rect 207900 42120 208000 42150
rect 204000 42100 204120 42120
rect 204380 42100 204620 42120
rect 204880 42100 205120 42120
rect 205380 42100 205620 42120
rect 205880 42100 206120 42120
rect 206380 42100 206620 42120
rect 206880 42100 207120 42120
rect 207380 42100 207620 42120
rect 207880 42100 208000 42120
rect 204000 42090 208000 42100
rect 204000 42020 204150 42090
rect 204350 42020 204650 42090
rect 204850 42020 205150 42090
rect 205350 42020 205650 42090
rect 205850 42020 206150 42090
rect 206350 42020 206650 42090
rect 206850 42020 207150 42090
rect 207350 42020 207650 42090
rect 207850 42020 208000 42090
rect 204000 41980 208000 42020
rect 204000 41910 204150 41980
rect 204350 41910 204650 41980
rect 204850 41910 205150 41980
rect 205350 41910 205650 41980
rect 205850 41910 206150 41980
rect 206350 41910 206650 41980
rect 206850 41910 207150 41980
rect 207350 41910 207650 41980
rect 207850 41910 208000 41980
rect 204000 41900 208000 41910
rect 204000 41880 204120 41900
rect 204380 41880 204620 41900
rect 204880 41880 205120 41900
rect 205380 41880 205620 41900
rect 205880 41880 206120 41900
rect 206380 41880 206620 41900
rect 206880 41880 207120 41900
rect 207380 41880 207620 41900
rect 207880 41880 208000 41900
rect 204000 41850 204100 41880
rect 204000 41650 204020 41850
rect 204090 41650 204100 41850
rect 204000 41620 204100 41650
rect 204400 41850 204600 41880
rect 204400 41650 204410 41850
rect 204480 41650 204520 41850
rect 204590 41650 204600 41850
rect 204400 41620 204600 41650
rect 204900 41850 205100 41880
rect 204900 41650 204910 41850
rect 204980 41650 205020 41850
rect 205090 41650 205100 41850
rect 204900 41620 205100 41650
rect 205400 41850 205600 41880
rect 205400 41650 205410 41850
rect 205480 41650 205520 41850
rect 205590 41650 205600 41850
rect 205400 41620 205600 41650
rect 205900 41850 206100 41880
rect 205900 41650 205910 41850
rect 205980 41650 206020 41850
rect 206090 41650 206100 41850
rect 205900 41620 206100 41650
rect 206400 41850 206600 41880
rect 206400 41650 206410 41850
rect 206480 41650 206520 41850
rect 206590 41650 206600 41850
rect 206400 41620 206600 41650
rect 206900 41850 207100 41880
rect 206900 41650 206910 41850
rect 206980 41650 207020 41850
rect 207090 41650 207100 41850
rect 206900 41620 207100 41650
rect 207400 41850 207600 41880
rect 207400 41650 207410 41850
rect 207480 41650 207520 41850
rect 207590 41650 207600 41850
rect 207400 41620 207600 41650
rect 207900 41850 208000 41880
rect 207900 41650 207910 41850
rect 207980 41650 208000 41850
rect 207900 41620 208000 41650
rect 204000 41600 204120 41620
rect 204380 41600 204620 41620
rect 204880 41600 205120 41620
rect 205380 41600 205620 41620
rect 205880 41600 206120 41620
rect 206380 41600 206620 41620
rect 206880 41600 207120 41620
rect 207380 41600 207620 41620
rect 207880 41600 208000 41620
rect 204000 41590 208000 41600
rect 204000 41520 204150 41590
rect 204350 41520 204650 41590
rect 204850 41520 205150 41590
rect 205350 41520 205650 41590
rect 205850 41520 206150 41590
rect 206350 41520 206650 41590
rect 206850 41520 207150 41590
rect 207350 41520 207650 41590
rect 207850 41520 208000 41590
rect 204000 41480 208000 41520
rect 204000 41410 204150 41480
rect 204350 41410 204650 41480
rect 204850 41410 205150 41480
rect 205350 41410 205650 41480
rect 205850 41410 206150 41480
rect 206350 41410 206650 41480
rect 206850 41410 207150 41480
rect 207350 41410 207650 41480
rect 207850 41410 208000 41480
rect 204000 41400 208000 41410
rect 204000 41380 204120 41400
rect 204380 41380 204620 41400
rect 204880 41380 205120 41400
rect 205380 41380 205620 41400
rect 205880 41380 206120 41400
rect 206380 41380 206620 41400
rect 206880 41380 207120 41400
rect 207380 41380 207620 41400
rect 207880 41380 208000 41400
rect 204000 41350 204100 41380
rect 204000 41150 204020 41350
rect 204090 41150 204100 41350
rect 204000 41120 204100 41150
rect 204400 41350 204600 41380
rect 204400 41150 204410 41350
rect 204480 41150 204520 41350
rect 204590 41150 204600 41350
rect 204400 41120 204600 41150
rect 204900 41350 205100 41380
rect 204900 41150 204910 41350
rect 204980 41150 205020 41350
rect 205090 41150 205100 41350
rect 204900 41120 205100 41150
rect 205400 41350 205600 41380
rect 205400 41150 205410 41350
rect 205480 41150 205520 41350
rect 205590 41150 205600 41350
rect 205400 41120 205600 41150
rect 205900 41350 206100 41380
rect 205900 41150 205910 41350
rect 205980 41150 206020 41350
rect 206090 41150 206100 41350
rect 205900 41120 206100 41150
rect 206400 41350 206600 41380
rect 206400 41150 206410 41350
rect 206480 41150 206520 41350
rect 206590 41150 206600 41350
rect 206400 41120 206600 41150
rect 206900 41350 207100 41380
rect 206900 41150 206910 41350
rect 206980 41150 207020 41350
rect 207090 41150 207100 41350
rect 206900 41120 207100 41150
rect 207400 41350 207600 41380
rect 207400 41150 207410 41350
rect 207480 41150 207520 41350
rect 207590 41150 207600 41350
rect 207400 41120 207600 41150
rect 207900 41350 208000 41380
rect 207900 41150 207910 41350
rect 207980 41150 208000 41350
rect 207900 41120 208000 41150
rect 204000 41100 204120 41120
rect 204380 41100 204620 41120
rect 204880 41100 205120 41120
rect 205380 41100 205620 41120
rect 205880 41100 206120 41120
rect 206380 41100 206620 41120
rect 206880 41100 207120 41120
rect 207380 41100 207620 41120
rect 207880 41100 208000 41120
rect 204000 41090 208000 41100
rect 204000 41020 204150 41090
rect 204350 41020 204650 41090
rect 204850 41020 205150 41090
rect 205350 41020 205650 41090
rect 205850 41020 206150 41090
rect 206350 41020 206650 41090
rect 206850 41020 207150 41090
rect 207350 41020 207650 41090
rect 207850 41020 208000 41090
rect 204000 40980 208000 41020
rect 204000 40910 204150 40980
rect 204350 40910 204650 40980
rect 204850 40910 205150 40980
rect 205350 40910 205650 40980
rect 205850 40910 206150 40980
rect 206350 40910 206650 40980
rect 206850 40910 207150 40980
rect 207350 40910 207650 40980
rect 207850 40910 208000 40980
rect 204000 40900 208000 40910
rect 204000 40880 204120 40900
rect 204380 40880 204620 40900
rect 204880 40880 205120 40900
rect 205380 40880 205620 40900
rect 205880 40880 206120 40900
rect 206380 40880 206620 40900
rect 206880 40880 207120 40900
rect 207380 40880 207620 40900
rect 207880 40880 208000 40900
rect 204000 40850 204100 40880
rect 204000 40650 204020 40850
rect 204090 40650 204100 40850
rect 204000 40620 204100 40650
rect 204400 40850 204600 40880
rect 204400 40650 204410 40850
rect 204480 40650 204520 40850
rect 204590 40650 204600 40850
rect 204400 40620 204600 40650
rect 204900 40850 205100 40880
rect 204900 40650 204910 40850
rect 204980 40650 205020 40850
rect 205090 40650 205100 40850
rect 204900 40620 205100 40650
rect 205400 40850 205600 40880
rect 205400 40650 205410 40850
rect 205480 40650 205520 40850
rect 205590 40650 205600 40850
rect 205400 40620 205600 40650
rect 205900 40850 206100 40880
rect 205900 40650 205910 40850
rect 205980 40650 206020 40850
rect 206090 40650 206100 40850
rect 205900 40620 206100 40650
rect 206400 40850 206600 40880
rect 206400 40650 206410 40850
rect 206480 40650 206520 40850
rect 206590 40650 206600 40850
rect 206400 40620 206600 40650
rect 206900 40850 207100 40880
rect 206900 40650 206910 40850
rect 206980 40650 207020 40850
rect 207090 40650 207100 40850
rect 206900 40620 207100 40650
rect 207400 40850 207600 40880
rect 207400 40650 207410 40850
rect 207480 40650 207520 40850
rect 207590 40650 207600 40850
rect 207400 40620 207600 40650
rect 207900 40850 208000 40880
rect 207900 40650 207910 40850
rect 207980 40650 208000 40850
rect 207900 40620 208000 40650
rect 204000 40600 204120 40620
rect 204380 40600 204620 40620
rect 204880 40600 205120 40620
rect 205380 40600 205620 40620
rect 205880 40600 206120 40620
rect 206380 40600 206620 40620
rect 206880 40600 207120 40620
rect 207380 40600 207620 40620
rect 207880 40600 208000 40620
rect 204000 40590 208000 40600
rect 204000 40520 204150 40590
rect 204350 40520 204650 40590
rect 204850 40520 205150 40590
rect 205350 40520 205650 40590
rect 205850 40520 206150 40590
rect 206350 40520 206650 40590
rect 206850 40520 207150 40590
rect 207350 40520 207650 40590
rect 207850 40520 208000 40590
rect 204000 40480 208000 40520
rect 204000 40410 204150 40480
rect 204350 40410 204650 40480
rect 204850 40410 205150 40480
rect 205350 40410 205650 40480
rect 205850 40410 206150 40480
rect 206350 40410 206650 40480
rect 206850 40410 207150 40480
rect 207350 40410 207650 40480
rect 207850 40410 208000 40480
rect 204000 40400 208000 40410
rect 204000 40380 204120 40400
rect 204380 40380 204620 40400
rect 204880 40380 205120 40400
rect 205380 40380 205620 40400
rect 205880 40380 206120 40400
rect 206380 40380 206620 40400
rect 206880 40380 207120 40400
rect 207380 40380 207620 40400
rect 207880 40380 208000 40400
rect 204000 40350 204100 40380
rect 204000 40150 204020 40350
rect 204090 40150 204100 40350
rect 204000 40120 204100 40150
rect 204400 40350 204600 40380
rect 204400 40150 204410 40350
rect 204480 40150 204520 40350
rect 204590 40150 204600 40350
rect 204400 40120 204600 40150
rect 204900 40350 205100 40380
rect 204900 40150 204910 40350
rect 204980 40150 205020 40350
rect 205090 40150 205100 40350
rect 204900 40120 205100 40150
rect 205400 40350 205600 40380
rect 205400 40150 205410 40350
rect 205480 40150 205520 40350
rect 205590 40150 205600 40350
rect 205400 40120 205600 40150
rect 205900 40350 206100 40380
rect 205900 40150 205910 40350
rect 205980 40150 206020 40350
rect 206090 40150 206100 40350
rect 205900 40120 206100 40150
rect 206400 40350 206600 40380
rect 206400 40150 206410 40350
rect 206480 40150 206520 40350
rect 206590 40150 206600 40350
rect 206400 40120 206600 40150
rect 206900 40350 207100 40380
rect 206900 40150 206910 40350
rect 206980 40150 207020 40350
rect 207090 40150 207100 40350
rect 206900 40120 207100 40150
rect 207400 40350 207600 40380
rect 207400 40150 207410 40350
rect 207480 40150 207520 40350
rect 207590 40150 207600 40350
rect 207400 40120 207600 40150
rect 207900 40350 208000 40380
rect 207900 40150 207910 40350
rect 207980 40150 208000 40350
rect 207900 40120 208000 40150
rect 204000 40100 204120 40120
rect 204380 40100 204620 40120
rect 204880 40100 205120 40120
rect 205380 40100 205620 40120
rect 205880 40100 206120 40120
rect 206380 40100 206620 40120
rect 206880 40100 207120 40120
rect 207380 40100 207620 40120
rect 207880 40100 208000 40120
rect 204000 40090 208000 40100
rect 204000 40020 204150 40090
rect 204350 40020 204650 40090
rect 204850 40020 205150 40090
rect 205350 40020 205650 40090
rect 205850 40020 206150 40090
rect 206350 40020 206650 40090
rect 206850 40020 207150 40090
rect 207350 40020 207650 40090
rect 207850 40020 208000 40090
rect 204000 39980 208000 40020
rect 204000 39910 204150 39980
rect 204350 39910 204650 39980
rect 204850 39910 205150 39980
rect 205350 39910 205650 39980
rect 205850 39910 206150 39980
rect 206350 39910 206650 39980
rect 206850 39910 207150 39980
rect 207350 39910 207650 39980
rect 207850 39910 208000 39980
rect 204000 39900 208000 39910
rect 204000 39880 204120 39900
rect 204380 39880 204620 39900
rect 204880 39880 205120 39900
rect 205380 39880 205620 39900
rect 205880 39880 206120 39900
rect 206380 39880 206620 39900
rect 206880 39880 207120 39900
rect 207380 39880 207620 39900
rect 207880 39880 208000 39900
rect 204000 39850 204100 39880
rect 204000 39650 204020 39850
rect 204090 39650 204100 39850
rect 204000 39620 204100 39650
rect 204400 39850 204600 39880
rect 204400 39650 204410 39850
rect 204480 39650 204520 39850
rect 204590 39650 204600 39850
rect 204400 39620 204600 39650
rect 204900 39850 205100 39880
rect 204900 39650 204910 39850
rect 204980 39650 205020 39850
rect 205090 39650 205100 39850
rect 204900 39620 205100 39650
rect 205400 39850 205600 39880
rect 205400 39650 205410 39850
rect 205480 39650 205520 39850
rect 205590 39650 205600 39850
rect 205400 39620 205600 39650
rect 205900 39850 206100 39880
rect 205900 39650 205910 39850
rect 205980 39650 206020 39850
rect 206090 39650 206100 39850
rect 205900 39620 206100 39650
rect 206400 39850 206600 39880
rect 206400 39650 206410 39850
rect 206480 39650 206520 39850
rect 206590 39650 206600 39850
rect 206400 39620 206600 39650
rect 206900 39850 207100 39880
rect 206900 39650 206910 39850
rect 206980 39650 207020 39850
rect 207090 39650 207100 39850
rect 206900 39620 207100 39650
rect 207400 39850 207600 39880
rect 207400 39650 207410 39850
rect 207480 39650 207520 39850
rect 207590 39650 207600 39850
rect 207400 39620 207600 39650
rect 207900 39850 208000 39880
rect 207900 39650 207910 39850
rect 207980 39650 208000 39850
rect 207900 39620 208000 39650
rect 204000 39600 204120 39620
rect 204380 39600 204620 39620
rect 204880 39600 205120 39620
rect 205380 39600 205620 39620
rect 205880 39600 206120 39620
rect 206380 39600 206620 39620
rect 206880 39600 207120 39620
rect 207380 39600 207620 39620
rect 207880 39600 208000 39620
rect 204000 39590 208000 39600
rect 204000 39520 204150 39590
rect 204350 39520 204650 39590
rect 204850 39520 205150 39590
rect 205350 39520 205650 39590
rect 205850 39520 206150 39590
rect 206350 39520 206650 39590
rect 206850 39520 207150 39590
rect 207350 39520 207650 39590
rect 207850 39520 208000 39590
rect 204000 39480 208000 39520
rect 204000 39410 204150 39480
rect 204350 39410 204650 39480
rect 204850 39410 205150 39480
rect 205350 39410 205650 39480
rect 205850 39410 206150 39480
rect 206350 39410 206650 39480
rect 206850 39410 207150 39480
rect 207350 39410 207650 39480
rect 207850 39410 208000 39480
rect 204000 39400 208000 39410
rect 204000 39380 204120 39400
rect 204380 39380 204620 39400
rect 204880 39380 205120 39400
rect 205380 39380 205620 39400
rect 205880 39380 206120 39400
rect 206380 39380 206620 39400
rect 206880 39380 207120 39400
rect 207380 39380 207620 39400
rect 207880 39380 208000 39400
rect 204000 39350 204100 39380
rect 204000 39150 204020 39350
rect 204090 39150 204100 39350
rect 204000 39120 204100 39150
rect 204400 39350 204600 39380
rect 204400 39150 204410 39350
rect 204480 39150 204520 39350
rect 204590 39150 204600 39350
rect 204400 39120 204600 39150
rect 204900 39350 205100 39380
rect 204900 39150 204910 39350
rect 204980 39150 205020 39350
rect 205090 39150 205100 39350
rect 204900 39120 205100 39150
rect 205400 39350 205600 39380
rect 205400 39150 205410 39350
rect 205480 39150 205520 39350
rect 205590 39150 205600 39350
rect 205400 39120 205600 39150
rect 205900 39350 206100 39380
rect 205900 39150 205910 39350
rect 205980 39150 206020 39350
rect 206090 39150 206100 39350
rect 205900 39120 206100 39150
rect 206400 39350 206600 39380
rect 206400 39150 206410 39350
rect 206480 39150 206520 39350
rect 206590 39150 206600 39350
rect 206400 39120 206600 39150
rect 206900 39350 207100 39380
rect 206900 39150 206910 39350
rect 206980 39150 207020 39350
rect 207090 39150 207100 39350
rect 206900 39120 207100 39150
rect 207400 39350 207600 39380
rect 207400 39150 207410 39350
rect 207480 39150 207520 39350
rect 207590 39150 207600 39350
rect 207400 39120 207600 39150
rect 207900 39350 208000 39380
rect 207900 39150 207910 39350
rect 207980 39150 208000 39350
rect 207900 39120 208000 39150
rect 204000 39100 204120 39120
rect 204380 39100 204620 39120
rect 204880 39100 205120 39120
rect 205380 39100 205620 39120
rect 205880 39100 206120 39120
rect 206380 39100 206620 39120
rect 206880 39100 207120 39120
rect 207380 39100 207620 39120
rect 207880 39100 208000 39120
rect 204000 39090 208000 39100
rect 204000 39020 204150 39090
rect 204350 39020 204650 39090
rect 204850 39020 205150 39090
rect 205350 39020 205650 39090
rect 205850 39020 206150 39090
rect 206350 39020 206650 39090
rect 206850 39020 207150 39090
rect 207350 39020 207650 39090
rect 207850 39020 208000 39090
rect 132000 38900 134000 39000
rect 132000 38880 132120 38900
rect 132380 38880 132620 38900
rect 132880 38880 133120 38900
rect 133380 38880 133620 38900
rect 133880 38880 134000 38900
rect 132000 38620 132100 38880
rect 132400 38620 132600 38880
rect 132900 38620 133100 38880
rect 133400 38620 133600 38880
rect 133900 38620 134000 38880
rect 132000 38600 132120 38620
rect 132380 38600 132620 38620
rect 132880 38600 133120 38620
rect 133380 38600 133620 38620
rect 133880 38600 134000 38620
rect 132000 38400 134000 38600
rect 132000 38380 132120 38400
rect 132380 38380 132620 38400
rect 132880 38380 133120 38400
rect 133380 38380 133620 38400
rect 133880 38380 134000 38400
rect 132000 38120 132100 38380
rect 132400 38120 132600 38380
rect 132900 38120 133100 38380
rect 133400 38120 133600 38380
rect 133900 38120 134000 38380
rect 132000 38100 132120 38120
rect 132380 38100 132620 38120
rect 132880 38100 133120 38120
rect 133380 38100 133620 38120
rect 133880 38100 134000 38120
rect 132000 37900 134000 38100
rect 132000 37880 132120 37900
rect 132380 37880 132620 37900
rect 132880 37880 133120 37900
rect 133380 37880 133620 37900
rect 133880 37880 134000 37900
rect 132000 37620 132100 37880
rect 132400 37620 132600 37880
rect 132900 37620 133100 37880
rect 133400 37620 133600 37880
rect 133900 37620 134000 37880
rect 132000 37600 132120 37620
rect 132380 37600 132620 37620
rect 132880 37600 133120 37620
rect 133380 37600 133620 37620
rect 133880 37600 134000 37620
rect 132000 37400 134000 37600
rect 132000 37380 132120 37400
rect 132380 37380 132620 37400
rect 132880 37380 133120 37400
rect 133380 37380 133620 37400
rect 133880 37380 134000 37400
rect 132000 37120 132100 37380
rect 132400 37120 132600 37380
rect 132900 37120 133100 37380
rect 133400 37120 133600 37380
rect 133900 37120 134000 37380
rect 132000 37100 132120 37120
rect 132380 37100 132620 37120
rect 132880 37100 133120 37120
rect 133380 37100 133620 37120
rect 133880 37100 134000 37120
rect 132000 36900 134000 37100
rect 132000 36880 132120 36900
rect 132380 36880 132620 36900
rect 132880 36880 133120 36900
rect 133380 36880 133620 36900
rect 133880 36880 134000 36900
rect 132000 36620 132100 36880
rect 132400 36620 132600 36880
rect 132900 36620 133100 36880
rect 133400 36620 133600 36880
rect 133900 36620 134000 36880
rect 132000 36600 132120 36620
rect 132380 36600 132620 36620
rect 132880 36600 133120 36620
rect 133380 36600 133620 36620
rect 133880 36600 134000 36620
rect 132000 36400 134000 36600
rect 132000 36380 132120 36400
rect 132380 36380 132620 36400
rect 132880 36380 133120 36400
rect 133380 36380 133620 36400
rect 133880 36380 134000 36400
rect 132000 36120 132100 36380
rect 132400 36120 132600 36380
rect 132900 36120 133100 36380
rect 133400 36120 133600 36380
rect 133900 36120 134000 36380
rect 132000 36100 132120 36120
rect 132380 36100 132620 36120
rect 132880 36100 133120 36120
rect 133380 36100 133620 36120
rect 133880 36100 134000 36120
rect 132000 35900 134000 36100
rect 132000 35880 132120 35900
rect 132380 35880 132620 35900
rect 132880 35880 133120 35900
rect 133380 35880 133620 35900
rect 133880 35880 134000 35900
rect 132000 35620 132100 35880
rect 132400 35620 132600 35880
rect 132900 35620 133100 35880
rect 133400 35620 133600 35880
rect 133900 35620 134000 35880
rect 132000 35600 132120 35620
rect 132380 35600 132620 35620
rect 132880 35600 133120 35620
rect 133380 35600 133620 35620
rect 133880 35600 134000 35620
rect 132000 35400 134000 35600
rect 132000 35380 132120 35400
rect 132380 35380 132620 35400
rect 132880 35380 133120 35400
rect 133380 35380 133620 35400
rect 133880 35380 134000 35400
rect 132000 35120 132100 35380
rect 132400 35120 132600 35380
rect 132900 35120 133100 35380
rect 133400 35120 133600 35380
rect 133900 35120 134000 35380
rect 132000 35100 132120 35120
rect 132380 35100 132620 35120
rect 132880 35100 133120 35120
rect 133380 35100 133620 35120
rect 133880 35100 134000 35120
rect 132000 34900 134000 35100
rect 132000 34880 132120 34900
rect 132380 34880 132620 34900
rect 132880 34880 133120 34900
rect 133380 34880 133620 34900
rect 133880 34880 134000 34900
rect 132000 34620 132100 34880
rect 132400 34620 132600 34880
rect 132900 34620 133100 34880
rect 133400 34620 133600 34880
rect 133900 34620 134000 34880
rect 132000 34600 132120 34620
rect 132380 34600 132620 34620
rect 132880 34600 133120 34620
rect 133380 34600 133620 34620
rect 133880 34600 134000 34620
rect 132000 34400 134000 34600
rect 132000 34380 132120 34400
rect 132380 34380 132620 34400
rect 132880 34380 133120 34400
rect 133380 34380 133620 34400
rect 133880 34380 134000 34400
rect 132000 34120 132100 34380
rect 132400 34120 132600 34380
rect 132900 34120 133100 34380
rect 133400 34120 133600 34380
rect 133900 34120 134000 34380
rect 132000 34100 132120 34120
rect 132380 34100 132620 34120
rect 132880 34100 133120 34120
rect 133380 34100 133620 34120
rect 133880 34100 134000 34120
rect 132000 33900 134000 34100
rect 132000 33880 132120 33900
rect 132380 33880 132620 33900
rect 132880 33880 133120 33900
rect 133380 33880 133620 33900
rect 133880 33880 134000 33900
rect 132000 33620 132100 33880
rect 132400 33620 132600 33880
rect 132900 33620 133100 33880
rect 133400 33620 133600 33880
rect 133900 33620 134000 33880
rect 132000 33600 132120 33620
rect 132380 33600 132620 33620
rect 132880 33600 133120 33620
rect 133380 33600 133620 33620
rect 133880 33600 134000 33620
rect 132000 33400 134000 33600
rect 132000 33380 132120 33400
rect 132380 33380 132620 33400
rect 132880 33380 133120 33400
rect 133380 33380 133620 33400
rect 133880 33380 134000 33400
rect 132000 33120 132100 33380
rect 132400 33120 132600 33380
rect 132900 33120 133100 33380
rect 133400 33120 133600 33380
rect 133900 33120 134000 33380
rect 132000 33100 132120 33120
rect 132380 33100 132620 33120
rect 132880 33100 133120 33120
rect 133380 33100 133620 33120
rect 133880 33100 134000 33120
rect 132000 33000 134000 33100
rect 204000 38980 208000 39020
rect 204000 38910 204150 38980
rect 204350 38910 204650 38980
rect 204850 38910 205150 38980
rect 205350 38910 205650 38980
rect 205850 38910 206150 38980
rect 206350 38910 206650 38980
rect 206850 38910 207150 38980
rect 207350 38910 207650 38980
rect 207850 38910 208000 38980
rect 204000 38900 208000 38910
rect 204000 38880 204120 38900
rect 204380 38880 204620 38900
rect 204880 38880 205120 38900
rect 205380 38880 205620 38900
rect 205880 38880 206120 38900
rect 206380 38880 206620 38900
rect 206880 38880 207120 38900
rect 207380 38880 207620 38900
rect 207880 38880 208000 38900
rect 204000 38850 204100 38880
rect 204000 38650 204020 38850
rect 204090 38650 204100 38850
rect 204000 38620 204100 38650
rect 204400 38850 204600 38880
rect 204400 38650 204410 38850
rect 204480 38650 204520 38850
rect 204590 38650 204600 38850
rect 204400 38620 204600 38650
rect 204900 38850 205100 38880
rect 204900 38650 204910 38850
rect 204980 38650 205020 38850
rect 205090 38650 205100 38850
rect 204900 38620 205100 38650
rect 205400 38850 205600 38880
rect 205400 38650 205410 38850
rect 205480 38650 205520 38850
rect 205590 38650 205600 38850
rect 205400 38620 205600 38650
rect 205900 38850 206100 38880
rect 205900 38650 205910 38850
rect 205980 38650 206020 38850
rect 206090 38650 206100 38850
rect 205900 38620 206100 38650
rect 206400 38850 206600 38880
rect 206400 38650 206410 38850
rect 206480 38650 206520 38850
rect 206590 38650 206600 38850
rect 206400 38620 206600 38650
rect 206900 38850 207100 38880
rect 206900 38650 206910 38850
rect 206980 38650 207020 38850
rect 207090 38650 207100 38850
rect 206900 38620 207100 38650
rect 207400 38850 207600 38880
rect 207400 38650 207410 38850
rect 207480 38650 207520 38850
rect 207590 38650 207600 38850
rect 207400 38620 207600 38650
rect 207900 38850 208000 38880
rect 207900 38650 207910 38850
rect 207980 38650 208000 38850
rect 207900 38620 208000 38650
rect 204000 38600 204120 38620
rect 204380 38600 204620 38620
rect 204880 38600 205120 38620
rect 205380 38600 205620 38620
rect 205880 38600 206120 38620
rect 206380 38600 206620 38620
rect 206880 38600 207120 38620
rect 207380 38600 207620 38620
rect 207880 38600 208000 38620
rect 204000 38590 208000 38600
rect 204000 38520 204150 38590
rect 204350 38520 204650 38590
rect 204850 38520 205150 38590
rect 205350 38520 205650 38590
rect 205850 38520 206150 38590
rect 206350 38520 206650 38590
rect 206850 38520 207150 38590
rect 207350 38520 207650 38590
rect 207850 38520 208000 38590
rect 204000 38480 208000 38520
rect 204000 38410 204150 38480
rect 204350 38410 204650 38480
rect 204850 38410 205150 38480
rect 205350 38410 205650 38480
rect 205850 38410 206150 38480
rect 206350 38410 206650 38480
rect 206850 38410 207150 38480
rect 207350 38410 207650 38480
rect 207850 38410 208000 38480
rect 204000 38400 208000 38410
rect 204000 38380 204120 38400
rect 204380 38380 204620 38400
rect 204880 38380 205120 38400
rect 205380 38380 205620 38400
rect 205880 38380 206120 38400
rect 206380 38380 206620 38400
rect 206880 38380 207120 38400
rect 207380 38380 207620 38400
rect 207880 38380 208000 38400
rect 204000 38350 204100 38380
rect 204000 38150 204020 38350
rect 204090 38150 204100 38350
rect 204000 38120 204100 38150
rect 204400 38350 204600 38380
rect 204400 38150 204410 38350
rect 204480 38150 204520 38350
rect 204590 38150 204600 38350
rect 204400 38120 204600 38150
rect 204900 38350 205100 38380
rect 204900 38150 204910 38350
rect 204980 38150 205020 38350
rect 205090 38150 205100 38350
rect 204900 38120 205100 38150
rect 205400 38350 205600 38380
rect 205400 38150 205410 38350
rect 205480 38150 205520 38350
rect 205590 38150 205600 38350
rect 205400 38120 205600 38150
rect 205900 38350 206100 38380
rect 205900 38150 205910 38350
rect 205980 38150 206020 38350
rect 206090 38150 206100 38350
rect 205900 38120 206100 38150
rect 206400 38350 206600 38380
rect 206400 38150 206410 38350
rect 206480 38150 206520 38350
rect 206590 38150 206600 38350
rect 206400 38120 206600 38150
rect 206900 38350 207100 38380
rect 206900 38150 206910 38350
rect 206980 38150 207020 38350
rect 207090 38150 207100 38350
rect 206900 38120 207100 38150
rect 207400 38350 207600 38380
rect 207400 38150 207410 38350
rect 207480 38150 207520 38350
rect 207590 38150 207600 38350
rect 207400 38120 207600 38150
rect 207900 38350 208000 38380
rect 207900 38150 207910 38350
rect 207980 38150 208000 38350
rect 207900 38120 208000 38150
rect 204000 38100 204120 38120
rect 204380 38100 204620 38120
rect 204880 38100 205120 38120
rect 205380 38100 205620 38120
rect 205880 38100 206120 38120
rect 206380 38100 206620 38120
rect 206880 38100 207120 38120
rect 207380 38100 207620 38120
rect 207880 38100 208000 38120
rect 204000 38090 208000 38100
rect 204000 38020 204150 38090
rect 204350 38020 204650 38090
rect 204850 38020 205150 38090
rect 205350 38020 205650 38090
rect 205850 38020 206150 38090
rect 206350 38020 206650 38090
rect 206850 38020 207150 38090
rect 207350 38020 207650 38090
rect 207850 38020 208000 38090
rect 204000 37980 208000 38020
rect 204000 37910 204150 37980
rect 204350 37910 204650 37980
rect 204850 37910 205150 37980
rect 205350 37910 205650 37980
rect 205850 37910 206150 37980
rect 206350 37910 206650 37980
rect 206850 37910 207150 37980
rect 207350 37910 207650 37980
rect 207850 37910 208000 37980
rect 204000 37900 208000 37910
rect 204000 37880 204120 37900
rect 204380 37880 204620 37900
rect 204880 37880 205120 37900
rect 205380 37880 205620 37900
rect 205880 37880 206120 37900
rect 206380 37880 206620 37900
rect 206880 37880 207120 37900
rect 207380 37880 207620 37900
rect 207880 37880 208000 37900
rect 204000 37850 204100 37880
rect 204000 37650 204020 37850
rect 204090 37650 204100 37850
rect 204000 37620 204100 37650
rect 204400 37850 204600 37880
rect 204400 37650 204410 37850
rect 204480 37650 204520 37850
rect 204590 37650 204600 37850
rect 204400 37620 204600 37650
rect 204900 37850 205100 37880
rect 204900 37650 204910 37850
rect 204980 37650 205020 37850
rect 205090 37650 205100 37850
rect 204900 37620 205100 37650
rect 205400 37850 205600 37880
rect 205400 37650 205410 37850
rect 205480 37650 205520 37850
rect 205590 37650 205600 37850
rect 205400 37620 205600 37650
rect 205900 37850 206100 37880
rect 205900 37650 205910 37850
rect 205980 37650 206020 37850
rect 206090 37650 206100 37850
rect 205900 37620 206100 37650
rect 206400 37850 206600 37880
rect 206400 37650 206410 37850
rect 206480 37650 206520 37850
rect 206590 37650 206600 37850
rect 206400 37620 206600 37650
rect 206900 37850 207100 37880
rect 206900 37650 206910 37850
rect 206980 37650 207020 37850
rect 207090 37650 207100 37850
rect 206900 37620 207100 37650
rect 207400 37850 207600 37880
rect 207400 37650 207410 37850
rect 207480 37650 207520 37850
rect 207590 37650 207600 37850
rect 207400 37620 207600 37650
rect 207900 37850 208000 37880
rect 207900 37650 207910 37850
rect 207980 37650 208000 37850
rect 207900 37620 208000 37650
rect 204000 37600 204120 37620
rect 204380 37600 204620 37620
rect 204880 37600 205120 37620
rect 205380 37600 205620 37620
rect 205880 37600 206120 37620
rect 206380 37600 206620 37620
rect 206880 37600 207120 37620
rect 207380 37600 207620 37620
rect 207880 37600 208000 37620
rect 204000 37590 208000 37600
rect 204000 37520 204150 37590
rect 204350 37520 204650 37590
rect 204850 37520 205150 37590
rect 205350 37520 205650 37590
rect 205850 37520 206150 37590
rect 206350 37520 206650 37590
rect 206850 37520 207150 37590
rect 207350 37520 207650 37590
rect 207850 37520 208000 37590
rect 204000 37480 208000 37520
rect 204000 37410 204150 37480
rect 204350 37410 204650 37480
rect 204850 37410 205150 37480
rect 205350 37410 205650 37480
rect 205850 37410 206150 37480
rect 206350 37410 206650 37480
rect 206850 37410 207150 37480
rect 207350 37410 207650 37480
rect 207850 37410 208000 37480
rect 204000 37400 208000 37410
rect 204000 37380 204120 37400
rect 204380 37380 204620 37400
rect 204880 37380 205120 37400
rect 205380 37380 205620 37400
rect 205880 37380 206120 37400
rect 206380 37380 206620 37400
rect 206880 37380 207120 37400
rect 207380 37380 207620 37400
rect 207880 37380 208000 37400
rect 204000 37350 204100 37380
rect 204000 37150 204020 37350
rect 204090 37150 204100 37350
rect 204000 37120 204100 37150
rect 204400 37350 204600 37380
rect 204400 37150 204410 37350
rect 204480 37150 204520 37350
rect 204590 37150 204600 37350
rect 204400 37120 204600 37150
rect 204900 37350 205100 37380
rect 204900 37150 204910 37350
rect 204980 37150 205020 37350
rect 205090 37150 205100 37350
rect 204900 37120 205100 37150
rect 205400 37350 205600 37380
rect 205400 37150 205410 37350
rect 205480 37150 205520 37350
rect 205590 37150 205600 37350
rect 205400 37120 205600 37150
rect 205900 37350 206100 37380
rect 205900 37150 205910 37350
rect 205980 37150 206020 37350
rect 206090 37150 206100 37350
rect 205900 37120 206100 37150
rect 206400 37350 206600 37380
rect 206400 37150 206410 37350
rect 206480 37150 206520 37350
rect 206590 37150 206600 37350
rect 206400 37120 206600 37150
rect 206900 37350 207100 37380
rect 206900 37150 206910 37350
rect 206980 37150 207020 37350
rect 207090 37150 207100 37350
rect 206900 37120 207100 37150
rect 207400 37350 207600 37380
rect 207400 37150 207410 37350
rect 207480 37150 207520 37350
rect 207590 37150 207600 37350
rect 207400 37120 207600 37150
rect 207900 37350 208000 37380
rect 207900 37150 207910 37350
rect 207980 37150 208000 37350
rect 207900 37120 208000 37150
rect 204000 37100 204120 37120
rect 204380 37100 204620 37120
rect 204880 37100 205120 37120
rect 205380 37100 205620 37120
rect 205880 37100 206120 37120
rect 206380 37100 206620 37120
rect 206880 37100 207120 37120
rect 207380 37100 207620 37120
rect 207880 37100 208000 37120
rect 204000 37090 208000 37100
rect 204000 37020 204150 37090
rect 204350 37020 204650 37090
rect 204850 37020 205150 37090
rect 205350 37020 205650 37090
rect 205850 37020 206150 37090
rect 206350 37020 206650 37090
rect 206850 37020 207150 37090
rect 207350 37020 207650 37090
rect 207850 37020 208000 37090
rect 204000 36980 208000 37020
rect 204000 36910 204150 36980
rect 204350 36910 204650 36980
rect 204850 36910 205150 36980
rect 205350 36910 205650 36980
rect 205850 36910 206150 36980
rect 206350 36910 206650 36980
rect 206850 36910 207150 36980
rect 207350 36910 207650 36980
rect 207850 36910 208000 36980
rect 204000 36900 208000 36910
rect 204000 36880 204120 36900
rect 204380 36880 204620 36900
rect 204880 36880 205120 36900
rect 205380 36880 205620 36900
rect 205880 36880 206120 36900
rect 206380 36880 206620 36900
rect 206880 36880 207120 36900
rect 207380 36880 207620 36900
rect 207880 36880 208000 36900
rect 204000 36850 204100 36880
rect 204000 36650 204020 36850
rect 204090 36650 204100 36850
rect 204000 36620 204100 36650
rect 204400 36850 204600 36880
rect 204400 36650 204410 36850
rect 204480 36650 204520 36850
rect 204590 36650 204600 36850
rect 204400 36620 204600 36650
rect 204900 36850 205100 36880
rect 204900 36650 204910 36850
rect 204980 36650 205020 36850
rect 205090 36650 205100 36850
rect 204900 36620 205100 36650
rect 205400 36850 205600 36880
rect 205400 36650 205410 36850
rect 205480 36650 205520 36850
rect 205590 36650 205600 36850
rect 205400 36620 205600 36650
rect 205900 36850 206100 36880
rect 205900 36650 205910 36850
rect 205980 36650 206020 36850
rect 206090 36650 206100 36850
rect 205900 36620 206100 36650
rect 206400 36850 206600 36880
rect 206400 36650 206410 36850
rect 206480 36650 206520 36850
rect 206590 36650 206600 36850
rect 206400 36620 206600 36650
rect 206900 36850 207100 36880
rect 206900 36650 206910 36850
rect 206980 36650 207020 36850
rect 207090 36650 207100 36850
rect 206900 36620 207100 36650
rect 207400 36850 207600 36880
rect 207400 36650 207410 36850
rect 207480 36650 207520 36850
rect 207590 36650 207600 36850
rect 207400 36620 207600 36650
rect 207900 36850 208000 36880
rect 207900 36650 207910 36850
rect 207980 36650 208000 36850
rect 207900 36620 208000 36650
rect 204000 36600 204120 36620
rect 204380 36600 204620 36620
rect 204880 36600 205120 36620
rect 205380 36600 205620 36620
rect 205880 36600 206120 36620
rect 206380 36600 206620 36620
rect 206880 36600 207120 36620
rect 207380 36600 207620 36620
rect 207880 36600 208000 36620
rect 204000 36590 208000 36600
rect 204000 36520 204150 36590
rect 204350 36520 204650 36590
rect 204850 36520 205150 36590
rect 205350 36520 205650 36590
rect 205850 36520 206150 36590
rect 206350 36520 206650 36590
rect 206850 36520 207150 36590
rect 207350 36520 207650 36590
rect 207850 36520 208000 36590
rect 204000 36480 208000 36520
rect 204000 36410 204150 36480
rect 204350 36410 204650 36480
rect 204850 36410 205150 36480
rect 205350 36410 205650 36480
rect 205850 36410 206150 36480
rect 206350 36410 206650 36480
rect 206850 36410 207150 36480
rect 207350 36410 207650 36480
rect 207850 36410 208000 36480
rect 204000 36400 208000 36410
rect 204000 36380 204120 36400
rect 204380 36380 204620 36400
rect 204880 36380 205120 36400
rect 205380 36380 205620 36400
rect 205880 36380 206120 36400
rect 206380 36380 206620 36400
rect 206880 36380 207120 36400
rect 207380 36380 207620 36400
rect 207880 36380 208000 36400
rect 204000 36350 204100 36380
rect 204000 36150 204020 36350
rect 204090 36150 204100 36350
rect 204000 36120 204100 36150
rect 204400 36350 204600 36380
rect 204400 36150 204410 36350
rect 204480 36150 204520 36350
rect 204590 36150 204600 36350
rect 204400 36120 204600 36150
rect 204900 36350 205100 36380
rect 204900 36150 204910 36350
rect 204980 36150 205020 36350
rect 205090 36150 205100 36350
rect 204900 36120 205100 36150
rect 205400 36350 205600 36380
rect 205400 36150 205410 36350
rect 205480 36150 205520 36350
rect 205590 36150 205600 36350
rect 205400 36120 205600 36150
rect 205900 36350 206100 36380
rect 205900 36150 205910 36350
rect 205980 36150 206020 36350
rect 206090 36150 206100 36350
rect 205900 36120 206100 36150
rect 206400 36350 206600 36380
rect 206400 36150 206410 36350
rect 206480 36150 206520 36350
rect 206590 36150 206600 36350
rect 206400 36120 206600 36150
rect 206900 36350 207100 36380
rect 206900 36150 206910 36350
rect 206980 36150 207020 36350
rect 207090 36150 207100 36350
rect 206900 36120 207100 36150
rect 207400 36350 207600 36380
rect 207400 36150 207410 36350
rect 207480 36150 207520 36350
rect 207590 36150 207600 36350
rect 207400 36120 207600 36150
rect 207900 36350 208000 36380
rect 207900 36150 207910 36350
rect 207980 36150 208000 36350
rect 207900 36120 208000 36150
rect 204000 36100 204120 36120
rect 204380 36100 204620 36120
rect 204880 36100 205120 36120
rect 205380 36100 205620 36120
rect 205880 36100 206120 36120
rect 206380 36100 206620 36120
rect 206880 36100 207120 36120
rect 207380 36100 207620 36120
rect 207880 36100 208000 36120
rect 204000 36090 208000 36100
rect 204000 36020 204150 36090
rect 204350 36020 204650 36090
rect 204850 36020 205150 36090
rect 205350 36020 205650 36090
rect 205850 36020 206150 36090
rect 206350 36020 206650 36090
rect 206850 36020 207150 36090
rect 207350 36020 207650 36090
rect 207850 36020 208000 36090
rect 204000 35980 208000 36020
rect 204000 35910 204150 35980
rect 204350 35910 204650 35980
rect 204850 35910 205150 35980
rect 205350 35910 205650 35980
rect 205850 35910 206150 35980
rect 206350 35910 206650 35980
rect 206850 35910 207150 35980
rect 207350 35910 207650 35980
rect 207850 35910 208000 35980
rect 204000 35900 208000 35910
rect 204000 35880 204120 35900
rect 204380 35880 204620 35900
rect 204880 35880 205120 35900
rect 205380 35880 205620 35900
rect 205880 35880 206120 35900
rect 206380 35880 206620 35900
rect 206880 35880 207120 35900
rect 207380 35880 207620 35900
rect 207880 35880 208000 35900
rect 204000 35850 204100 35880
rect 204000 35650 204020 35850
rect 204090 35650 204100 35850
rect 204000 35620 204100 35650
rect 204400 35850 204600 35880
rect 204400 35650 204410 35850
rect 204480 35650 204520 35850
rect 204590 35650 204600 35850
rect 204400 35620 204600 35650
rect 204900 35850 205100 35880
rect 204900 35650 204910 35850
rect 204980 35650 205020 35850
rect 205090 35650 205100 35850
rect 204900 35620 205100 35650
rect 205400 35850 205600 35880
rect 205400 35650 205410 35850
rect 205480 35650 205520 35850
rect 205590 35650 205600 35850
rect 205400 35620 205600 35650
rect 205900 35850 206100 35880
rect 205900 35650 205910 35850
rect 205980 35650 206020 35850
rect 206090 35650 206100 35850
rect 205900 35620 206100 35650
rect 206400 35850 206600 35880
rect 206400 35650 206410 35850
rect 206480 35650 206520 35850
rect 206590 35650 206600 35850
rect 206400 35620 206600 35650
rect 206900 35850 207100 35880
rect 206900 35650 206910 35850
rect 206980 35650 207020 35850
rect 207090 35650 207100 35850
rect 206900 35620 207100 35650
rect 207400 35850 207600 35880
rect 207400 35650 207410 35850
rect 207480 35650 207520 35850
rect 207590 35650 207600 35850
rect 207400 35620 207600 35650
rect 207900 35850 208000 35880
rect 207900 35650 207910 35850
rect 207980 35650 208000 35850
rect 207900 35620 208000 35650
rect 204000 35600 204120 35620
rect 204380 35600 204620 35620
rect 204880 35600 205120 35620
rect 205380 35600 205620 35620
rect 205880 35600 206120 35620
rect 206380 35600 206620 35620
rect 206880 35600 207120 35620
rect 207380 35600 207620 35620
rect 207880 35600 208000 35620
rect 204000 35590 208000 35600
rect 204000 35520 204150 35590
rect 204350 35520 204650 35590
rect 204850 35520 205150 35590
rect 205350 35520 205650 35590
rect 205850 35520 206150 35590
rect 206350 35520 206650 35590
rect 206850 35520 207150 35590
rect 207350 35520 207650 35590
rect 207850 35520 208000 35590
rect 204000 35480 208000 35520
rect 204000 35410 204150 35480
rect 204350 35410 204650 35480
rect 204850 35410 205150 35480
rect 205350 35410 205650 35480
rect 205850 35410 206150 35480
rect 206350 35410 206650 35480
rect 206850 35410 207150 35480
rect 207350 35410 207650 35480
rect 207850 35410 208000 35480
rect 204000 35400 208000 35410
rect 204000 35380 204120 35400
rect 204380 35380 204620 35400
rect 204880 35380 205120 35400
rect 205380 35380 205620 35400
rect 205880 35380 206120 35400
rect 206380 35380 206620 35400
rect 206880 35380 207120 35400
rect 207380 35380 207620 35400
rect 207880 35380 208000 35400
rect 204000 35350 204100 35380
rect 204000 35150 204020 35350
rect 204090 35150 204100 35350
rect 204000 35120 204100 35150
rect 204400 35350 204600 35380
rect 204400 35150 204410 35350
rect 204480 35150 204520 35350
rect 204590 35150 204600 35350
rect 204400 35120 204600 35150
rect 204900 35350 205100 35380
rect 204900 35150 204910 35350
rect 204980 35150 205020 35350
rect 205090 35150 205100 35350
rect 204900 35120 205100 35150
rect 205400 35350 205600 35380
rect 205400 35150 205410 35350
rect 205480 35150 205520 35350
rect 205590 35150 205600 35350
rect 205400 35120 205600 35150
rect 205900 35350 206100 35380
rect 205900 35150 205910 35350
rect 205980 35150 206020 35350
rect 206090 35150 206100 35350
rect 205900 35120 206100 35150
rect 206400 35350 206600 35380
rect 206400 35150 206410 35350
rect 206480 35150 206520 35350
rect 206590 35150 206600 35350
rect 206400 35120 206600 35150
rect 206900 35350 207100 35380
rect 206900 35150 206910 35350
rect 206980 35150 207020 35350
rect 207090 35150 207100 35350
rect 206900 35120 207100 35150
rect 207400 35350 207600 35380
rect 207400 35150 207410 35350
rect 207480 35150 207520 35350
rect 207590 35150 207600 35350
rect 207400 35120 207600 35150
rect 207900 35350 208000 35380
rect 207900 35150 207910 35350
rect 207980 35150 208000 35350
rect 207900 35120 208000 35150
rect 204000 35100 204120 35120
rect 204380 35100 204620 35120
rect 204880 35100 205120 35120
rect 205380 35100 205620 35120
rect 205880 35100 206120 35120
rect 206380 35100 206620 35120
rect 206880 35100 207120 35120
rect 207380 35100 207620 35120
rect 207880 35100 208000 35120
rect 204000 35090 208000 35100
rect 204000 35020 204150 35090
rect 204350 35020 204650 35090
rect 204850 35020 205150 35090
rect 205350 35020 205650 35090
rect 205850 35020 206150 35090
rect 206350 35020 206650 35090
rect 206850 35020 207150 35090
rect 207350 35020 207650 35090
rect 207850 35020 208000 35090
rect 204000 34980 208000 35020
rect 204000 34910 204150 34980
rect 204350 34910 204650 34980
rect 204850 34910 205150 34980
rect 205350 34910 205650 34980
rect 205850 34910 206150 34980
rect 206350 34910 206650 34980
rect 206850 34910 207150 34980
rect 207350 34910 207650 34980
rect 207850 34910 208000 34980
rect 204000 34900 208000 34910
rect 204000 34880 204120 34900
rect 204380 34880 204620 34900
rect 204880 34880 205120 34900
rect 205380 34880 205620 34900
rect 205880 34880 206120 34900
rect 206380 34880 206620 34900
rect 206880 34880 207120 34900
rect 207380 34880 207620 34900
rect 207880 34880 208000 34900
rect 204000 34850 204100 34880
rect 204000 34650 204020 34850
rect 204090 34650 204100 34850
rect 204000 34620 204100 34650
rect 204400 34850 204600 34880
rect 204400 34650 204410 34850
rect 204480 34650 204520 34850
rect 204590 34650 204600 34850
rect 204400 34620 204600 34650
rect 204900 34850 205100 34880
rect 204900 34650 204910 34850
rect 204980 34650 205020 34850
rect 205090 34650 205100 34850
rect 204900 34620 205100 34650
rect 205400 34850 205600 34880
rect 205400 34650 205410 34850
rect 205480 34650 205520 34850
rect 205590 34650 205600 34850
rect 205400 34620 205600 34650
rect 205900 34850 206100 34880
rect 205900 34650 205910 34850
rect 205980 34650 206020 34850
rect 206090 34650 206100 34850
rect 205900 34620 206100 34650
rect 206400 34850 206600 34880
rect 206400 34650 206410 34850
rect 206480 34650 206520 34850
rect 206590 34650 206600 34850
rect 206400 34620 206600 34650
rect 206900 34850 207100 34880
rect 206900 34650 206910 34850
rect 206980 34650 207020 34850
rect 207090 34650 207100 34850
rect 206900 34620 207100 34650
rect 207400 34850 207600 34880
rect 207400 34650 207410 34850
rect 207480 34650 207520 34850
rect 207590 34650 207600 34850
rect 207400 34620 207600 34650
rect 207900 34850 208000 34880
rect 207900 34650 207910 34850
rect 207980 34650 208000 34850
rect 207900 34620 208000 34650
rect 204000 34600 204120 34620
rect 204380 34600 204620 34620
rect 204880 34600 205120 34620
rect 205380 34600 205620 34620
rect 205880 34600 206120 34620
rect 206380 34600 206620 34620
rect 206880 34600 207120 34620
rect 207380 34600 207620 34620
rect 207880 34600 208000 34620
rect 204000 34590 208000 34600
rect 204000 34520 204150 34590
rect 204350 34520 204650 34590
rect 204850 34520 205150 34590
rect 205350 34520 205650 34590
rect 205850 34520 206150 34590
rect 206350 34520 206650 34590
rect 206850 34520 207150 34590
rect 207350 34520 207650 34590
rect 207850 34520 208000 34590
rect 204000 34480 208000 34520
rect 204000 34410 204150 34480
rect 204350 34410 204650 34480
rect 204850 34410 205150 34480
rect 205350 34410 205650 34480
rect 205850 34410 206150 34480
rect 206350 34410 206650 34480
rect 206850 34410 207150 34480
rect 207350 34410 207650 34480
rect 207850 34410 208000 34480
rect 204000 34400 208000 34410
rect 204000 34380 204120 34400
rect 204380 34380 204620 34400
rect 204880 34380 205120 34400
rect 205380 34380 205620 34400
rect 205880 34380 206120 34400
rect 206380 34380 206620 34400
rect 206880 34380 207120 34400
rect 207380 34380 207620 34400
rect 207880 34380 208000 34400
rect 204000 34350 204100 34380
rect 204000 34150 204020 34350
rect 204090 34150 204100 34350
rect 204000 34120 204100 34150
rect 204400 34350 204600 34380
rect 204400 34150 204410 34350
rect 204480 34150 204520 34350
rect 204590 34150 204600 34350
rect 204400 34120 204600 34150
rect 204900 34350 205100 34380
rect 204900 34150 204910 34350
rect 204980 34150 205020 34350
rect 205090 34150 205100 34350
rect 204900 34120 205100 34150
rect 205400 34350 205600 34380
rect 205400 34150 205410 34350
rect 205480 34150 205520 34350
rect 205590 34150 205600 34350
rect 205400 34120 205600 34150
rect 205900 34350 206100 34380
rect 205900 34150 205910 34350
rect 205980 34150 206020 34350
rect 206090 34150 206100 34350
rect 205900 34120 206100 34150
rect 206400 34350 206600 34380
rect 206400 34150 206410 34350
rect 206480 34150 206520 34350
rect 206590 34150 206600 34350
rect 206400 34120 206600 34150
rect 206900 34350 207100 34380
rect 206900 34150 206910 34350
rect 206980 34150 207020 34350
rect 207090 34150 207100 34350
rect 206900 34120 207100 34150
rect 207400 34350 207600 34380
rect 207400 34150 207410 34350
rect 207480 34150 207520 34350
rect 207590 34150 207600 34350
rect 207400 34120 207600 34150
rect 207900 34350 208000 34380
rect 207900 34150 207910 34350
rect 207980 34150 208000 34350
rect 207900 34120 208000 34150
rect 204000 34100 204120 34120
rect 204380 34100 204620 34120
rect 204880 34100 205120 34120
rect 205380 34100 205620 34120
rect 205880 34100 206120 34120
rect 206380 34100 206620 34120
rect 206880 34100 207120 34120
rect 207380 34100 207620 34120
rect 207880 34100 208000 34120
rect 204000 34090 208000 34100
rect 204000 34020 204150 34090
rect 204350 34020 204650 34090
rect 204850 34020 205150 34090
rect 205350 34020 205650 34090
rect 205850 34020 206150 34090
rect 206350 34020 206650 34090
rect 206850 34020 207150 34090
rect 207350 34020 207650 34090
rect 207850 34020 208000 34090
rect 204000 33980 208000 34020
rect 204000 33910 204150 33980
rect 204350 33910 204650 33980
rect 204850 33910 205150 33980
rect 205350 33910 205650 33980
rect 205850 33910 206150 33980
rect 206350 33910 206650 33980
rect 206850 33910 207150 33980
rect 207350 33910 207650 33980
rect 207850 33910 208000 33980
rect 204000 33900 208000 33910
rect 204000 33880 204120 33900
rect 204380 33880 204620 33900
rect 204880 33880 205120 33900
rect 205380 33880 205620 33900
rect 205880 33880 206120 33900
rect 206380 33880 206620 33900
rect 206880 33880 207120 33900
rect 207380 33880 207620 33900
rect 207880 33880 208000 33900
rect 204000 33850 204100 33880
rect 204000 33650 204020 33850
rect 204090 33650 204100 33850
rect 204000 33620 204100 33650
rect 204400 33850 204600 33880
rect 204400 33650 204410 33850
rect 204480 33650 204520 33850
rect 204590 33650 204600 33850
rect 204400 33620 204600 33650
rect 204900 33850 205100 33880
rect 204900 33650 204910 33850
rect 204980 33650 205020 33850
rect 205090 33650 205100 33850
rect 204900 33620 205100 33650
rect 205400 33850 205600 33880
rect 205400 33650 205410 33850
rect 205480 33650 205520 33850
rect 205590 33650 205600 33850
rect 205400 33620 205600 33650
rect 205900 33850 206100 33880
rect 205900 33650 205910 33850
rect 205980 33650 206020 33850
rect 206090 33650 206100 33850
rect 205900 33620 206100 33650
rect 206400 33850 206600 33880
rect 206400 33650 206410 33850
rect 206480 33650 206520 33850
rect 206590 33650 206600 33850
rect 206400 33620 206600 33650
rect 206900 33850 207100 33880
rect 206900 33650 206910 33850
rect 206980 33650 207020 33850
rect 207090 33650 207100 33850
rect 206900 33620 207100 33650
rect 207400 33850 207600 33880
rect 207400 33650 207410 33850
rect 207480 33650 207520 33850
rect 207590 33650 207600 33850
rect 207400 33620 207600 33650
rect 207900 33850 208000 33880
rect 207900 33650 207910 33850
rect 207980 33650 208000 33850
rect 207900 33620 208000 33650
rect 204000 33600 204120 33620
rect 204380 33600 204620 33620
rect 204880 33600 205120 33620
rect 205380 33600 205620 33620
rect 205880 33600 206120 33620
rect 206380 33600 206620 33620
rect 206880 33600 207120 33620
rect 207380 33600 207620 33620
rect 207880 33600 208000 33620
rect 204000 33590 208000 33600
rect 204000 33520 204150 33590
rect 204350 33520 204650 33590
rect 204850 33520 205150 33590
rect 205350 33520 205650 33590
rect 205850 33520 206150 33590
rect 206350 33520 206650 33590
rect 206850 33520 207150 33590
rect 207350 33520 207650 33590
rect 207850 33520 208000 33590
rect 204000 33480 208000 33520
rect 204000 33410 204150 33480
rect 204350 33410 204650 33480
rect 204850 33410 205150 33480
rect 205350 33410 205650 33480
rect 205850 33410 206150 33480
rect 206350 33410 206650 33480
rect 206850 33410 207150 33480
rect 207350 33410 207650 33480
rect 207850 33410 208000 33480
rect 204000 33400 208000 33410
rect 204000 33380 204120 33400
rect 204380 33380 204620 33400
rect 204880 33380 205120 33400
rect 205380 33380 205620 33400
rect 205880 33380 206120 33400
rect 206380 33380 206620 33400
rect 206880 33380 207120 33400
rect 207380 33380 207620 33400
rect 207880 33380 208000 33400
rect 204000 33350 204100 33380
rect 204000 33150 204020 33350
rect 204090 33150 204100 33350
rect 204000 33120 204100 33150
rect 204400 33350 204600 33380
rect 204400 33150 204410 33350
rect 204480 33150 204520 33350
rect 204590 33150 204600 33350
rect 204400 33120 204600 33150
rect 204900 33350 205100 33380
rect 204900 33150 204910 33350
rect 204980 33150 205020 33350
rect 205090 33150 205100 33350
rect 204900 33120 205100 33150
rect 205400 33350 205600 33380
rect 205400 33150 205410 33350
rect 205480 33150 205520 33350
rect 205590 33150 205600 33350
rect 205400 33120 205600 33150
rect 205900 33350 206100 33380
rect 205900 33150 205910 33350
rect 205980 33150 206020 33350
rect 206090 33150 206100 33350
rect 205900 33120 206100 33150
rect 206400 33350 206600 33380
rect 206400 33150 206410 33350
rect 206480 33150 206520 33350
rect 206590 33150 206600 33350
rect 206400 33120 206600 33150
rect 206900 33350 207100 33380
rect 206900 33150 206910 33350
rect 206980 33150 207020 33350
rect 207090 33150 207100 33350
rect 206900 33120 207100 33150
rect 207400 33350 207600 33380
rect 207400 33150 207410 33350
rect 207480 33150 207520 33350
rect 207590 33150 207600 33350
rect 207400 33120 207600 33150
rect 207900 33350 208000 33380
rect 207900 33150 207910 33350
rect 207980 33150 208000 33350
rect 207900 33120 208000 33150
rect 204000 33100 204120 33120
rect 204380 33100 204620 33120
rect 204880 33100 205120 33120
rect 205380 33100 205620 33120
rect 205880 33100 206120 33120
rect 206380 33100 206620 33120
rect 206880 33100 207120 33120
rect 207380 33100 207620 33120
rect 207880 33100 208000 33120
rect 204000 33090 208000 33100
rect 204000 33020 204150 33090
rect 204350 33020 204650 33090
rect 204850 33020 205150 33090
rect 205350 33020 205650 33090
rect 205850 33020 206150 33090
rect 206350 33020 206650 33090
rect 206850 33020 207150 33090
rect 207350 33020 207650 33090
rect 207850 33020 208000 33090
rect 132000 32900 138000 33000
rect 132000 32880 132120 32900
rect 132380 32880 132620 32900
rect 132880 32880 133120 32900
rect 133380 32880 133620 32900
rect 133880 32880 134120 32900
rect 134380 32880 134620 32900
rect 134880 32880 135120 32900
rect 135380 32880 135620 32900
rect 135880 32880 136120 32900
rect 136380 32880 136620 32900
rect 136880 32880 137120 32900
rect 137380 32880 137620 32900
rect 137880 32880 138000 32900
rect 132000 32620 132100 32880
rect 132400 32620 132600 32880
rect 132900 32620 133100 32880
rect 133400 32620 133600 32880
rect 133900 32620 134100 32880
rect 134400 32620 134600 32880
rect 134900 32620 135100 32880
rect 135400 32620 135600 32880
rect 135900 32620 136100 32880
rect 136400 32620 136600 32880
rect 136900 32620 137100 32880
rect 137400 32620 137600 32880
rect 137900 32620 138000 32880
rect 132000 32600 132120 32620
rect 132380 32600 132620 32620
rect 132880 32600 133120 32620
rect 133380 32600 133620 32620
rect 133880 32600 134120 32620
rect 134380 32600 134620 32620
rect 134880 32600 135120 32620
rect 135380 32600 135620 32620
rect 135880 32600 136120 32620
rect 136380 32600 136620 32620
rect 136880 32600 137120 32620
rect 137380 32600 137620 32620
rect 137880 32600 138000 32620
rect 132000 32400 138000 32600
rect 132000 32380 132120 32400
rect 132380 32380 132620 32400
rect 132880 32380 133120 32400
rect 133380 32380 133620 32400
rect 133880 32380 134120 32400
rect 134380 32380 134620 32400
rect 134880 32380 135120 32400
rect 135380 32380 135620 32400
rect 135880 32380 136120 32400
rect 136380 32380 136620 32400
rect 136880 32380 137120 32400
rect 137380 32380 137620 32400
rect 137880 32380 138000 32400
rect 132000 32120 132100 32380
rect 132400 32120 132600 32380
rect 132900 32120 133100 32380
rect 133400 32120 133600 32380
rect 133900 32120 134100 32380
rect 134400 32120 134600 32380
rect 134900 32120 135100 32380
rect 135400 32120 135600 32380
rect 135900 32120 136100 32380
rect 136400 32120 136600 32380
rect 136900 32120 137100 32380
rect 137400 32120 137600 32380
rect 137900 32120 138000 32380
rect 132000 32100 132120 32120
rect 132380 32100 132620 32120
rect 132880 32100 133120 32120
rect 133380 32100 133620 32120
rect 133880 32100 134120 32120
rect 134380 32100 134620 32120
rect 134880 32100 135120 32120
rect 135380 32100 135620 32120
rect 135880 32100 136120 32120
rect 136380 32100 136620 32120
rect 136880 32100 137120 32120
rect 137380 32100 137620 32120
rect 137880 32100 138000 32120
rect 132000 32000 138000 32100
rect 204000 32980 208000 33020
rect 204000 32910 204150 32980
rect 204350 32910 204650 32980
rect 204850 32910 205150 32980
rect 205350 32910 205650 32980
rect 205850 32910 206150 32980
rect 206350 32910 206650 32980
rect 206850 32910 207150 32980
rect 207350 32910 207650 32980
rect 207850 32910 208000 32980
rect 204000 32900 208000 32910
rect 204000 32880 204120 32900
rect 204380 32880 204620 32900
rect 204880 32880 205120 32900
rect 205380 32880 205620 32900
rect 205880 32880 206120 32900
rect 206380 32880 206620 32900
rect 206880 32880 207120 32900
rect 207380 32880 207620 32900
rect 207880 32880 208000 32900
rect 204000 32850 204100 32880
rect 204000 32650 204020 32850
rect 204090 32650 204100 32850
rect 204000 32620 204100 32650
rect 204400 32850 204600 32880
rect 204400 32650 204410 32850
rect 204480 32650 204520 32850
rect 204590 32650 204600 32850
rect 204400 32620 204600 32650
rect 204900 32850 205100 32880
rect 204900 32650 204910 32850
rect 204980 32650 205020 32850
rect 205090 32650 205100 32850
rect 204900 32620 205100 32650
rect 205400 32850 205600 32880
rect 205400 32650 205410 32850
rect 205480 32650 205520 32850
rect 205590 32650 205600 32850
rect 205400 32620 205600 32650
rect 205900 32850 206100 32880
rect 205900 32650 205910 32850
rect 205980 32650 206020 32850
rect 206090 32650 206100 32850
rect 205900 32620 206100 32650
rect 206400 32850 206600 32880
rect 206400 32650 206410 32850
rect 206480 32650 206520 32850
rect 206590 32650 206600 32850
rect 206400 32620 206600 32650
rect 206900 32850 207100 32880
rect 206900 32650 206910 32850
rect 206980 32650 207020 32850
rect 207090 32650 207100 32850
rect 206900 32620 207100 32650
rect 207400 32850 207600 32880
rect 207400 32650 207410 32850
rect 207480 32650 207520 32850
rect 207590 32650 207600 32850
rect 207400 32620 207600 32650
rect 207900 32850 208000 32880
rect 207900 32650 207910 32850
rect 207980 32650 208000 32850
rect 207900 32620 208000 32650
rect 204000 32600 204120 32620
rect 204380 32600 204620 32620
rect 204880 32600 205120 32620
rect 205380 32600 205620 32620
rect 205880 32600 206120 32620
rect 206380 32600 206620 32620
rect 206880 32600 207120 32620
rect 207380 32600 207620 32620
rect 207880 32600 208000 32620
rect 204000 32590 208000 32600
rect 204000 32520 204150 32590
rect 204350 32520 204650 32590
rect 204850 32520 205150 32590
rect 205350 32520 205650 32590
rect 205850 32520 206150 32590
rect 206350 32520 206650 32590
rect 206850 32520 207150 32590
rect 207350 32520 207650 32590
rect 207850 32520 208000 32590
rect 204000 32480 208000 32520
rect 204000 32410 204150 32480
rect 204350 32410 204650 32480
rect 204850 32410 205150 32480
rect 205350 32410 205650 32480
rect 205850 32410 206150 32480
rect 206350 32410 206650 32480
rect 206850 32410 207150 32480
rect 207350 32410 207650 32480
rect 207850 32410 208000 32480
rect 204000 32400 208000 32410
rect 204000 32380 204120 32400
rect 204380 32380 204620 32400
rect 204880 32380 205120 32400
rect 205380 32380 205620 32400
rect 205880 32380 206120 32400
rect 206380 32380 206620 32400
rect 206880 32380 207120 32400
rect 207380 32380 207620 32400
rect 207880 32380 208000 32400
rect 204000 32350 204100 32380
rect 204000 32150 204020 32350
rect 204090 32150 204100 32350
rect 204000 32120 204100 32150
rect 204400 32350 204600 32380
rect 204400 32150 204410 32350
rect 204480 32150 204520 32350
rect 204590 32150 204600 32350
rect 204400 32120 204600 32150
rect 204900 32350 205100 32380
rect 204900 32150 204910 32350
rect 204980 32150 205020 32350
rect 205090 32150 205100 32350
rect 204900 32120 205100 32150
rect 205400 32350 205600 32380
rect 205400 32150 205410 32350
rect 205480 32150 205520 32350
rect 205590 32150 205600 32350
rect 205400 32120 205600 32150
rect 205900 32350 206100 32380
rect 205900 32150 205910 32350
rect 205980 32150 206020 32350
rect 206090 32150 206100 32350
rect 205900 32120 206100 32150
rect 206400 32350 206600 32380
rect 206400 32150 206410 32350
rect 206480 32150 206520 32350
rect 206590 32150 206600 32350
rect 206400 32120 206600 32150
rect 206900 32350 207100 32380
rect 206900 32150 206910 32350
rect 206980 32150 207020 32350
rect 207090 32150 207100 32350
rect 206900 32120 207100 32150
rect 207400 32350 207600 32380
rect 207400 32150 207410 32350
rect 207480 32150 207520 32350
rect 207590 32150 207600 32350
rect 207400 32120 207600 32150
rect 207900 32350 208000 32380
rect 207900 32150 207910 32350
rect 207980 32150 208000 32350
rect 207900 32120 208000 32150
rect 204000 32100 204120 32120
rect 204380 32100 204620 32120
rect 204880 32100 205120 32120
rect 205380 32100 205620 32120
rect 205880 32100 206120 32120
rect 206380 32100 206620 32120
rect 206880 32100 207120 32120
rect 207380 32100 207620 32120
rect 207880 32100 208000 32120
rect 204000 32090 208000 32100
rect 204000 32020 204150 32090
rect 204350 32020 204650 32090
rect 204850 32020 205150 32090
rect 205350 32020 205650 32090
rect 205850 32020 206150 32090
rect 206350 32020 206650 32090
rect 206850 32020 207150 32090
rect 207350 32020 207650 32090
rect 207850 32020 208000 32090
rect 134000 31900 140000 32000
rect 134000 31880 134120 31900
rect 134380 31880 134620 31900
rect 134880 31880 135120 31900
rect 135380 31880 135620 31900
rect 135880 31880 136120 31900
rect 136380 31880 136620 31900
rect 136880 31880 137120 31900
rect 137380 31880 137620 31900
rect 137880 31880 138120 31900
rect 138380 31880 138620 31900
rect 138880 31880 139120 31900
rect 139380 31880 139620 31900
rect 139880 31880 140000 31900
rect 134000 31620 134100 31880
rect 134400 31620 134600 31880
rect 134900 31620 135100 31880
rect 135400 31620 135600 31880
rect 135900 31620 136100 31880
rect 136400 31620 136600 31880
rect 136900 31620 137100 31880
rect 137400 31620 137600 31880
rect 137900 31620 138100 31880
rect 138400 31620 138600 31880
rect 138900 31620 139100 31880
rect 139400 31620 139600 31880
rect 139900 31620 140000 31880
rect 134000 31600 134120 31620
rect 134380 31600 134620 31620
rect 134880 31600 135120 31620
rect 135380 31600 135620 31620
rect 135880 31600 136120 31620
rect 136380 31600 136620 31620
rect 136880 31600 137120 31620
rect 137380 31600 137620 31620
rect 137880 31600 138120 31620
rect 138380 31600 138620 31620
rect 138880 31600 139120 31620
rect 139380 31600 139620 31620
rect 139880 31600 140000 31620
rect 134000 31400 140000 31600
rect 134000 31380 134120 31400
rect 134380 31380 134620 31400
rect 134880 31380 135120 31400
rect 135380 31380 135620 31400
rect 135880 31380 136120 31400
rect 136380 31380 136620 31400
rect 136880 31380 137120 31400
rect 137380 31380 137620 31400
rect 137880 31380 138120 31400
rect 138380 31380 138620 31400
rect 138880 31380 139120 31400
rect 139380 31380 139620 31400
rect 139880 31380 140000 31400
rect 134000 31120 134100 31380
rect 134400 31120 134600 31380
rect 134900 31120 135100 31380
rect 135400 31120 135600 31380
rect 135900 31120 136100 31380
rect 136400 31120 136600 31380
rect 136900 31120 137100 31380
rect 137400 31120 137600 31380
rect 137900 31120 138100 31380
rect 138400 31120 138600 31380
rect 138900 31120 139100 31380
rect 139400 31120 139600 31380
rect 139900 31120 140000 31380
rect 134000 31100 134120 31120
rect 134380 31100 134620 31120
rect 134880 31100 135120 31120
rect 135380 31100 135620 31120
rect 135880 31100 136120 31120
rect 136380 31100 136620 31120
rect 136880 31100 137120 31120
rect 137380 31100 137620 31120
rect 137880 31100 138120 31120
rect 138380 31100 138620 31120
rect 138880 31100 139120 31120
rect 139380 31100 139620 31120
rect 139880 31100 140000 31120
rect 134000 30900 140000 31100
rect 134000 30880 134120 30900
rect 134380 30880 134620 30900
rect 134880 30880 135120 30900
rect 135380 30880 135620 30900
rect 135880 30880 136120 30900
rect 136380 30880 136620 30900
rect 136880 30880 137120 30900
rect 137380 30880 137620 30900
rect 137880 30880 138120 30900
rect 138380 30880 138620 30900
rect 138880 30880 139120 30900
rect 139380 30880 139620 30900
rect 139880 30880 140000 30900
rect 134000 30620 134100 30880
rect 134400 30620 134600 30880
rect 134900 30620 135100 30880
rect 135400 30620 135600 30880
rect 135900 30620 136100 30880
rect 136400 30620 136600 30880
rect 136900 30620 137100 30880
rect 137400 30620 137600 30880
rect 137900 30620 138100 30880
rect 138400 30620 138600 30880
rect 138900 30620 139100 30880
rect 139400 30620 139600 30880
rect 139900 30620 140000 30880
rect 134000 30600 134120 30620
rect 134380 30600 134620 30620
rect 134880 30600 135120 30620
rect 135380 30600 135620 30620
rect 135880 30600 136120 30620
rect 136380 30600 136620 30620
rect 136880 30600 137120 30620
rect 137380 30600 137620 30620
rect 137880 30600 138120 30620
rect 138380 30600 138620 30620
rect 138880 30600 139120 30620
rect 139380 30600 139620 30620
rect 139880 30600 140000 30620
rect 134000 30400 140000 30600
rect 134000 30380 134120 30400
rect 134380 30380 134620 30400
rect 134880 30380 135120 30400
rect 135380 30380 135620 30400
rect 135880 30380 136120 30400
rect 136380 30380 136620 30400
rect 136880 30380 137120 30400
rect 137380 30380 137620 30400
rect 137880 30380 138120 30400
rect 138380 30380 138620 30400
rect 138880 30380 139120 30400
rect 139380 30380 139620 30400
rect 139880 30380 140000 30400
rect 134000 30120 134100 30380
rect 134400 30120 134600 30380
rect 134900 30120 135100 30380
rect 135400 30120 135600 30380
rect 135900 30120 136100 30380
rect 136400 30120 136600 30380
rect 136900 30120 137100 30380
rect 137400 30120 137600 30380
rect 137900 30120 138100 30380
rect 138400 30120 138600 30380
rect 138900 30120 139100 30380
rect 139400 30120 139600 30380
rect 139900 30120 140000 30380
rect 134000 30100 134120 30120
rect 134380 30100 134620 30120
rect 134880 30100 135120 30120
rect 135380 30100 135620 30120
rect 135880 30100 136120 30120
rect 136380 30100 136620 30120
rect 136880 30100 137120 30120
rect 137380 30100 137620 30120
rect 137880 30100 138120 30120
rect 138380 30100 138620 30120
rect 138880 30100 139120 30120
rect 139380 30100 139620 30120
rect 139880 30100 140000 30120
rect 134000 30000 140000 30100
rect 204000 31980 208000 32020
rect 204000 31910 204150 31980
rect 204350 31910 204650 31980
rect 204850 31910 205150 31980
rect 205350 31910 205650 31980
rect 205850 31910 206150 31980
rect 206350 31910 206650 31980
rect 206850 31910 207150 31980
rect 207350 31910 207650 31980
rect 207850 31910 208000 31980
rect 204000 31900 208000 31910
rect 204000 31880 204120 31900
rect 204380 31880 204620 31900
rect 204880 31880 205120 31900
rect 205380 31880 205620 31900
rect 205880 31880 206120 31900
rect 206380 31880 206620 31900
rect 206880 31880 207120 31900
rect 207380 31880 207620 31900
rect 207880 31880 208000 31900
rect 204000 31850 204100 31880
rect 204000 31650 204020 31850
rect 204090 31650 204100 31850
rect 204000 31620 204100 31650
rect 204400 31850 204600 31880
rect 204400 31650 204410 31850
rect 204480 31650 204520 31850
rect 204590 31650 204600 31850
rect 204400 31620 204600 31650
rect 204900 31850 205100 31880
rect 204900 31650 204910 31850
rect 204980 31650 205020 31850
rect 205090 31650 205100 31850
rect 204900 31620 205100 31650
rect 205400 31850 205600 31880
rect 205400 31650 205410 31850
rect 205480 31650 205520 31850
rect 205590 31650 205600 31850
rect 205400 31620 205600 31650
rect 205900 31850 206100 31880
rect 205900 31650 205910 31850
rect 205980 31650 206020 31850
rect 206090 31650 206100 31850
rect 205900 31620 206100 31650
rect 206400 31850 206600 31880
rect 206400 31650 206410 31850
rect 206480 31650 206520 31850
rect 206590 31650 206600 31850
rect 206400 31620 206600 31650
rect 206900 31850 207100 31880
rect 206900 31650 206910 31850
rect 206980 31650 207020 31850
rect 207090 31650 207100 31850
rect 206900 31620 207100 31650
rect 207400 31850 207600 31880
rect 207400 31650 207410 31850
rect 207480 31650 207520 31850
rect 207590 31650 207600 31850
rect 207400 31620 207600 31650
rect 207900 31850 208000 31880
rect 207900 31650 207910 31850
rect 207980 31650 208000 31850
rect 207900 31620 208000 31650
rect 204000 31600 204120 31620
rect 204380 31600 204620 31620
rect 204880 31600 205120 31620
rect 205380 31600 205620 31620
rect 205880 31600 206120 31620
rect 206380 31600 206620 31620
rect 206880 31600 207120 31620
rect 207380 31600 207620 31620
rect 207880 31600 208000 31620
rect 204000 31590 208000 31600
rect 204000 31520 204150 31590
rect 204350 31520 204650 31590
rect 204850 31520 205150 31590
rect 205350 31520 205650 31590
rect 205850 31520 206150 31590
rect 206350 31520 206650 31590
rect 206850 31520 207150 31590
rect 207350 31520 207650 31590
rect 207850 31520 208000 31590
rect 204000 31480 208000 31520
rect 204000 31410 204150 31480
rect 204350 31410 204650 31480
rect 204850 31410 205150 31480
rect 205350 31410 205650 31480
rect 205850 31410 206150 31480
rect 206350 31410 206650 31480
rect 206850 31410 207150 31480
rect 207350 31410 207650 31480
rect 207850 31410 208000 31480
rect 204000 31400 208000 31410
rect 204000 31380 204120 31400
rect 204380 31380 204620 31400
rect 204880 31380 205120 31400
rect 205380 31380 205620 31400
rect 205880 31380 206120 31400
rect 206380 31380 206620 31400
rect 206880 31380 207120 31400
rect 207380 31380 207620 31400
rect 207880 31380 208000 31400
rect 204000 31350 204100 31380
rect 204000 31150 204020 31350
rect 204090 31150 204100 31350
rect 204000 31120 204100 31150
rect 204400 31350 204600 31380
rect 204400 31150 204410 31350
rect 204480 31150 204520 31350
rect 204590 31150 204600 31350
rect 204400 31120 204600 31150
rect 204900 31350 205100 31380
rect 204900 31150 204910 31350
rect 204980 31150 205020 31350
rect 205090 31150 205100 31350
rect 204900 31120 205100 31150
rect 205400 31350 205600 31380
rect 205400 31150 205410 31350
rect 205480 31150 205520 31350
rect 205590 31150 205600 31350
rect 205400 31120 205600 31150
rect 205900 31350 206100 31380
rect 205900 31150 205910 31350
rect 205980 31150 206020 31350
rect 206090 31150 206100 31350
rect 205900 31120 206100 31150
rect 206400 31350 206600 31380
rect 206400 31150 206410 31350
rect 206480 31150 206520 31350
rect 206590 31150 206600 31350
rect 206400 31120 206600 31150
rect 206900 31350 207100 31380
rect 206900 31150 206910 31350
rect 206980 31150 207020 31350
rect 207090 31150 207100 31350
rect 206900 31120 207100 31150
rect 207400 31350 207600 31380
rect 207400 31150 207410 31350
rect 207480 31150 207520 31350
rect 207590 31150 207600 31350
rect 207400 31120 207600 31150
rect 207900 31350 208000 31380
rect 207900 31150 207910 31350
rect 207980 31150 208000 31350
rect 207900 31120 208000 31150
rect 204000 31100 204120 31120
rect 204380 31100 204620 31120
rect 204880 31100 205120 31120
rect 205380 31100 205620 31120
rect 205880 31100 206120 31120
rect 206380 31100 206620 31120
rect 206880 31100 207120 31120
rect 207380 31100 207620 31120
rect 207880 31100 208000 31120
rect 204000 31090 208000 31100
rect 204000 31020 204150 31090
rect 204350 31020 204650 31090
rect 204850 31020 205150 31090
rect 205350 31020 205650 31090
rect 205850 31020 206150 31090
rect 206350 31020 206650 31090
rect 206850 31020 207150 31090
rect 207350 31020 207650 31090
rect 207850 31020 208000 31090
rect 204000 30980 208000 31020
rect 204000 30910 204150 30980
rect 204350 30910 204650 30980
rect 204850 30910 205150 30980
rect 205350 30910 205650 30980
rect 205850 30910 206150 30980
rect 206350 30910 206650 30980
rect 206850 30910 207150 30980
rect 207350 30910 207650 30980
rect 207850 30910 208000 30980
rect 204000 30900 208000 30910
rect 204000 30880 204120 30900
rect 204380 30880 204620 30900
rect 204880 30880 205120 30900
rect 205380 30880 205620 30900
rect 205880 30880 206120 30900
rect 206380 30880 206620 30900
rect 206880 30880 207120 30900
rect 207380 30880 207620 30900
rect 207880 30880 208000 30900
rect 204000 30850 204100 30880
rect 204000 30650 204020 30850
rect 204090 30650 204100 30850
rect 204000 30620 204100 30650
rect 204400 30850 204600 30880
rect 204400 30650 204410 30850
rect 204480 30650 204520 30850
rect 204590 30650 204600 30850
rect 204400 30620 204600 30650
rect 204900 30850 205100 30880
rect 204900 30650 204910 30850
rect 204980 30650 205020 30850
rect 205090 30650 205100 30850
rect 204900 30620 205100 30650
rect 205400 30850 205600 30880
rect 205400 30650 205410 30850
rect 205480 30650 205520 30850
rect 205590 30650 205600 30850
rect 205400 30620 205600 30650
rect 205900 30850 206100 30880
rect 205900 30650 205910 30850
rect 205980 30650 206020 30850
rect 206090 30650 206100 30850
rect 205900 30620 206100 30650
rect 206400 30850 206600 30880
rect 206400 30650 206410 30850
rect 206480 30650 206520 30850
rect 206590 30650 206600 30850
rect 206400 30620 206600 30650
rect 206900 30850 207100 30880
rect 206900 30650 206910 30850
rect 206980 30650 207020 30850
rect 207090 30650 207100 30850
rect 206900 30620 207100 30650
rect 207400 30850 207600 30880
rect 207400 30650 207410 30850
rect 207480 30650 207520 30850
rect 207590 30650 207600 30850
rect 207400 30620 207600 30650
rect 207900 30850 208000 30880
rect 207900 30650 207910 30850
rect 207980 30650 208000 30850
rect 207900 30620 208000 30650
rect 204000 30600 204120 30620
rect 204380 30600 204620 30620
rect 204880 30600 205120 30620
rect 205380 30600 205620 30620
rect 205880 30600 206120 30620
rect 206380 30600 206620 30620
rect 206880 30600 207120 30620
rect 207380 30600 207620 30620
rect 207880 30600 208000 30620
rect 204000 30590 208000 30600
rect 204000 30520 204150 30590
rect 204350 30520 204650 30590
rect 204850 30520 205150 30590
rect 205350 30520 205650 30590
rect 205850 30520 206150 30590
rect 206350 30520 206650 30590
rect 206850 30520 207150 30590
rect 207350 30520 207650 30590
rect 207850 30520 208000 30590
rect 204000 30480 208000 30520
rect 204000 30410 204150 30480
rect 204350 30410 204650 30480
rect 204850 30410 205150 30480
rect 205350 30410 205650 30480
rect 205850 30410 206150 30480
rect 206350 30410 206650 30480
rect 206850 30410 207150 30480
rect 207350 30410 207650 30480
rect 207850 30410 208000 30480
rect 204000 30400 208000 30410
rect 204000 30380 204120 30400
rect 204380 30380 204620 30400
rect 204880 30380 205120 30400
rect 205380 30380 205620 30400
rect 205880 30380 206120 30400
rect 206380 30380 206620 30400
rect 206880 30380 207120 30400
rect 207380 30380 207620 30400
rect 207880 30380 208000 30400
rect 204000 30350 204100 30380
rect 204000 30150 204020 30350
rect 204090 30150 204100 30350
rect 204000 30120 204100 30150
rect 204400 30350 204600 30380
rect 204400 30150 204410 30350
rect 204480 30150 204520 30350
rect 204590 30150 204600 30350
rect 204400 30120 204600 30150
rect 204900 30350 205100 30380
rect 204900 30150 204910 30350
rect 204980 30150 205020 30350
rect 205090 30150 205100 30350
rect 204900 30120 205100 30150
rect 205400 30350 205600 30380
rect 205400 30150 205410 30350
rect 205480 30150 205520 30350
rect 205590 30150 205600 30350
rect 205400 30120 205600 30150
rect 205900 30350 206100 30380
rect 205900 30150 205910 30350
rect 205980 30150 206020 30350
rect 206090 30150 206100 30350
rect 205900 30120 206100 30150
rect 206400 30350 206600 30380
rect 206400 30150 206410 30350
rect 206480 30150 206520 30350
rect 206590 30150 206600 30350
rect 206400 30120 206600 30150
rect 206900 30350 207100 30380
rect 206900 30150 206910 30350
rect 206980 30150 207020 30350
rect 207090 30150 207100 30350
rect 206900 30120 207100 30150
rect 207400 30350 207600 30380
rect 207400 30150 207410 30350
rect 207480 30150 207520 30350
rect 207590 30150 207600 30350
rect 207400 30120 207600 30150
rect 207900 30350 208000 30380
rect 207900 30150 207910 30350
rect 207980 30150 208000 30350
rect 207900 30120 208000 30150
rect 204000 30100 204120 30120
rect 204380 30100 204620 30120
rect 204880 30100 205120 30120
rect 205380 30100 205620 30120
rect 205880 30100 206120 30120
rect 206380 30100 206620 30120
rect 206880 30100 207120 30120
rect 207380 30100 207620 30120
rect 207880 30100 208000 30120
rect 204000 30090 208000 30100
rect 204000 30020 204150 30090
rect 204350 30020 204650 30090
rect 204850 30020 205150 30090
rect 205350 30020 205650 30090
rect 205850 30020 206150 30090
rect 206350 30020 206650 30090
rect 206850 30020 207150 30090
rect 207350 30020 207650 30090
rect 207850 30020 208000 30090
rect 204000 29980 208000 30020
rect 204000 29910 204150 29980
rect 204350 29910 204650 29980
rect 204850 29910 205150 29980
rect 205350 29910 205650 29980
rect 205850 29910 206150 29980
rect 206350 29910 206650 29980
rect 206850 29910 207150 29980
rect 207350 29910 207650 29980
rect 207850 29910 208000 29980
rect 204000 29900 208000 29910
rect 204000 29880 204120 29900
rect 204380 29880 204620 29900
rect 204880 29880 205120 29900
rect 205380 29880 205620 29900
rect 205880 29880 206120 29900
rect 206380 29880 206620 29900
rect 206880 29880 207120 29900
rect 207380 29880 207620 29900
rect 207880 29880 208000 29900
rect 204000 29850 204100 29880
rect 204000 29650 204020 29850
rect 204090 29650 204100 29850
rect 204000 29620 204100 29650
rect 204400 29850 204600 29880
rect 204400 29650 204410 29850
rect 204480 29650 204520 29850
rect 204590 29650 204600 29850
rect 204400 29620 204600 29650
rect 204900 29850 205100 29880
rect 204900 29650 204910 29850
rect 204980 29650 205020 29850
rect 205090 29650 205100 29850
rect 204900 29620 205100 29650
rect 205400 29850 205600 29880
rect 205400 29650 205410 29850
rect 205480 29650 205520 29850
rect 205590 29650 205600 29850
rect 205400 29620 205600 29650
rect 205900 29850 206100 29880
rect 205900 29650 205910 29850
rect 205980 29650 206020 29850
rect 206090 29650 206100 29850
rect 205900 29620 206100 29650
rect 206400 29850 206600 29880
rect 206400 29650 206410 29850
rect 206480 29650 206520 29850
rect 206590 29650 206600 29850
rect 206400 29620 206600 29650
rect 206900 29850 207100 29880
rect 206900 29650 206910 29850
rect 206980 29650 207020 29850
rect 207090 29650 207100 29850
rect 206900 29620 207100 29650
rect 207400 29850 207600 29880
rect 207400 29650 207410 29850
rect 207480 29650 207520 29850
rect 207590 29650 207600 29850
rect 207400 29620 207600 29650
rect 207900 29850 208000 29880
rect 207900 29650 207910 29850
rect 207980 29650 208000 29850
rect 207900 29620 208000 29650
rect 204000 29600 204120 29620
rect 204380 29600 204620 29620
rect 204880 29600 205120 29620
rect 205380 29600 205620 29620
rect 205880 29600 206120 29620
rect 206380 29600 206620 29620
rect 206880 29600 207120 29620
rect 207380 29600 207620 29620
rect 207880 29600 208000 29620
rect 204000 29590 208000 29600
rect 204000 29520 204150 29590
rect 204350 29520 204650 29590
rect 204850 29520 205150 29590
rect 205350 29520 205650 29590
rect 205850 29520 206150 29590
rect 206350 29520 206650 29590
rect 206850 29520 207150 29590
rect 207350 29520 207650 29590
rect 207850 29520 208000 29590
rect 204000 29480 208000 29520
rect 204000 29410 204150 29480
rect 204350 29410 204650 29480
rect 204850 29410 205150 29480
rect 205350 29410 205650 29480
rect 205850 29410 206150 29480
rect 206350 29410 206650 29480
rect 206850 29410 207150 29480
rect 207350 29410 207650 29480
rect 207850 29410 208000 29480
rect 204000 29400 208000 29410
rect 204000 29380 204120 29400
rect 204380 29380 204620 29400
rect 204880 29380 205120 29400
rect 205380 29380 205620 29400
rect 205880 29380 206120 29400
rect 206380 29380 206620 29400
rect 206880 29380 207120 29400
rect 207380 29380 207620 29400
rect 207880 29380 208000 29400
rect 204000 29350 204100 29380
rect 204000 29150 204020 29350
rect 204090 29150 204100 29350
rect 204000 29120 204100 29150
rect 204400 29350 204600 29380
rect 204400 29150 204410 29350
rect 204480 29150 204520 29350
rect 204590 29150 204600 29350
rect 204400 29120 204600 29150
rect 204900 29350 205100 29380
rect 204900 29150 204910 29350
rect 204980 29150 205020 29350
rect 205090 29150 205100 29350
rect 204900 29120 205100 29150
rect 205400 29350 205600 29380
rect 205400 29150 205410 29350
rect 205480 29150 205520 29350
rect 205590 29150 205600 29350
rect 205400 29120 205600 29150
rect 205900 29350 206100 29380
rect 205900 29150 205910 29350
rect 205980 29150 206020 29350
rect 206090 29150 206100 29350
rect 205900 29120 206100 29150
rect 206400 29350 206600 29380
rect 206400 29150 206410 29350
rect 206480 29150 206520 29350
rect 206590 29150 206600 29350
rect 206400 29120 206600 29150
rect 206900 29350 207100 29380
rect 206900 29150 206910 29350
rect 206980 29150 207020 29350
rect 207090 29150 207100 29350
rect 206900 29120 207100 29150
rect 207400 29350 207600 29380
rect 207400 29150 207410 29350
rect 207480 29150 207520 29350
rect 207590 29150 207600 29350
rect 207400 29120 207600 29150
rect 207900 29350 208000 29380
rect 207900 29150 207910 29350
rect 207980 29150 208000 29350
rect 207900 29120 208000 29150
rect 204000 29100 204120 29120
rect 204380 29100 204620 29120
rect 204880 29100 205120 29120
rect 205380 29100 205620 29120
rect 205880 29100 206120 29120
rect 206380 29100 206620 29120
rect 206880 29100 207120 29120
rect 207380 29100 207620 29120
rect 207880 29100 208000 29120
rect 204000 29090 208000 29100
rect 204000 29020 204150 29090
rect 204350 29020 204650 29090
rect 204850 29020 205150 29090
rect 205350 29020 205650 29090
rect 205850 29020 206150 29090
rect 206350 29020 206650 29090
rect 206850 29020 207150 29090
rect 207350 29020 207650 29090
rect 207850 29020 208000 29090
rect 204000 28980 208000 29020
rect 204000 28910 204150 28980
rect 204350 28910 204650 28980
rect 204850 28910 205150 28980
rect 205350 28910 205650 28980
rect 205850 28910 206150 28980
rect 206350 28910 206650 28980
rect 206850 28910 207150 28980
rect 207350 28910 207650 28980
rect 207850 28910 208000 28980
rect 204000 28900 208000 28910
rect 204000 28880 204120 28900
rect 204380 28880 204620 28900
rect 204880 28880 205120 28900
rect 205380 28880 205620 28900
rect 205880 28880 206120 28900
rect 206380 28880 206620 28900
rect 206880 28880 207120 28900
rect 207380 28880 207620 28900
rect 207880 28880 208000 28900
rect 204000 28850 204100 28880
rect 204000 28650 204020 28850
rect 204090 28650 204100 28850
rect 204000 28620 204100 28650
rect 204400 28850 204600 28880
rect 204400 28650 204410 28850
rect 204480 28650 204520 28850
rect 204590 28650 204600 28850
rect 204400 28620 204600 28650
rect 204900 28850 205100 28880
rect 204900 28650 204910 28850
rect 204980 28650 205020 28850
rect 205090 28650 205100 28850
rect 204900 28620 205100 28650
rect 205400 28850 205600 28880
rect 205400 28650 205410 28850
rect 205480 28650 205520 28850
rect 205590 28650 205600 28850
rect 205400 28620 205600 28650
rect 205900 28850 206100 28880
rect 205900 28650 205910 28850
rect 205980 28650 206020 28850
rect 206090 28650 206100 28850
rect 205900 28620 206100 28650
rect 206400 28850 206600 28880
rect 206400 28650 206410 28850
rect 206480 28650 206520 28850
rect 206590 28650 206600 28850
rect 206400 28620 206600 28650
rect 206900 28850 207100 28880
rect 206900 28650 206910 28850
rect 206980 28650 207020 28850
rect 207090 28650 207100 28850
rect 206900 28620 207100 28650
rect 207400 28850 207600 28880
rect 207400 28650 207410 28850
rect 207480 28650 207520 28850
rect 207590 28650 207600 28850
rect 207400 28620 207600 28650
rect 207900 28850 208000 28880
rect 207900 28650 207910 28850
rect 207980 28650 208000 28850
rect 207900 28620 208000 28650
rect 204000 28600 204120 28620
rect 204380 28600 204620 28620
rect 204880 28600 205120 28620
rect 205380 28600 205620 28620
rect 205880 28600 206120 28620
rect 206380 28600 206620 28620
rect 206880 28600 207120 28620
rect 207380 28600 207620 28620
rect 207880 28600 208000 28620
rect 204000 28590 208000 28600
rect 204000 28520 204150 28590
rect 204350 28520 204650 28590
rect 204850 28520 205150 28590
rect 205350 28520 205650 28590
rect 205850 28520 206150 28590
rect 206350 28520 206650 28590
rect 206850 28520 207150 28590
rect 207350 28520 207650 28590
rect 207850 28520 208000 28590
rect 204000 28480 208000 28520
rect 204000 28410 204150 28480
rect 204350 28410 204650 28480
rect 204850 28410 205150 28480
rect 205350 28410 205650 28480
rect 205850 28410 206150 28480
rect 206350 28410 206650 28480
rect 206850 28410 207150 28480
rect 207350 28410 207650 28480
rect 207850 28410 208000 28480
rect 204000 28400 208000 28410
rect 204000 28380 204120 28400
rect 204380 28380 204620 28400
rect 204880 28380 205120 28400
rect 205380 28380 205620 28400
rect 205880 28380 206120 28400
rect 206380 28380 206620 28400
rect 206880 28380 207120 28400
rect 207380 28380 207620 28400
rect 207880 28380 208000 28400
rect 204000 28350 204100 28380
rect 204000 28150 204020 28350
rect 204090 28150 204100 28350
rect 204000 28120 204100 28150
rect 204400 28350 204600 28380
rect 204400 28150 204410 28350
rect 204480 28150 204520 28350
rect 204590 28150 204600 28350
rect 204400 28120 204600 28150
rect 204900 28350 205100 28380
rect 204900 28150 204910 28350
rect 204980 28150 205020 28350
rect 205090 28150 205100 28350
rect 204900 28120 205100 28150
rect 205400 28350 205600 28380
rect 205400 28150 205410 28350
rect 205480 28150 205520 28350
rect 205590 28150 205600 28350
rect 205400 28120 205600 28150
rect 205900 28350 206100 28380
rect 205900 28150 205910 28350
rect 205980 28150 206020 28350
rect 206090 28150 206100 28350
rect 205900 28120 206100 28150
rect 206400 28350 206600 28380
rect 206400 28150 206410 28350
rect 206480 28150 206520 28350
rect 206590 28150 206600 28350
rect 206400 28120 206600 28150
rect 206900 28350 207100 28380
rect 206900 28150 206910 28350
rect 206980 28150 207020 28350
rect 207090 28150 207100 28350
rect 206900 28120 207100 28150
rect 207400 28350 207600 28380
rect 207400 28150 207410 28350
rect 207480 28150 207520 28350
rect 207590 28150 207600 28350
rect 207400 28120 207600 28150
rect 207900 28350 208000 28380
rect 207900 28150 207910 28350
rect 207980 28150 208000 28350
rect 207900 28120 208000 28150
rect 204000 28100 204120 28120
rect 204380 28100 204620 28120
rect 204880 28100 205120 28120
rect 205380 28100 205620 28120
rect 205880 28100 206120 28120
rect 206380 28100 206620 28120
rect 206880 28100 207120 28120
rect 207380 28100 207620 28120
rect 207880 28100 208000 28120
rect 204000 28090 208000 28100
rect 204000 28020 204150 28090
rect 204350 28020 204650 28090
rect 204850 28020 205150 28090
rect 205350 28020 205650 28090
rect 205850 28020 206150 28090
rect 206350 28020 206650 28090
rect 206850 28020 207150 28090
rect 207350 28020 207650 28090
rect 207850 28020 208000 28090
rect 204000 27980 208000 28020
rect 204000 27910 204150 27980
rect 204350 27910 204650 27980
rect 204850 27910 205150 27980
rect 205350 27910 205650 27980
rect 205850 27910 206150 27980
rect 206350 27910 206650 27980
rect 206850 27910 207150 27980
rect 207350 27910 207650 27980
rect 207850 27910 208000 27980
rect 204000 27900 208000 27910
rect 204000 27880 204120 27900
rect 204380 27880 204620 27900
rect 204880 27880 205120 27900
rect 205380 27880 205620 27900
rect 205880 27880 206120 27900
rect 206380 27880 206620 27900
rect 206880 27880 207120 27900
rect 207380 27880 207620 27900
rect 207880 27880 208000 27900
rect 204000 27850 204100 27880
rect 204000 27650 204020 27850
rect 204090 27650 204100 27850
rect 204000 27620 204100 27650
rect 204400 27850 204600 27880
rect 204400 27650 204410 27850
rect 204480 27650 204520 27850
rect 204590 27650 204600 27850
rect 204400 27620 204600 27650
rect 204900 27850 205100 27880
rect 204900 27650 204910 27850
rect 204980 27650 205020 27850
rect 205090 27650 205100 27850
rect 204900 27620 205100 27650
rect 205400 27850 205600 27880
rect 205400 27650 205410 27850
rect 205480 27650 205520 27850
rect 205590 27650 205600 27850
rect 205400 27620 205600 27650
rect 205900 27850 206100 27880
rect 205900 27650 205910 27850
rect 205980 27650 206020 27850
rect 206090 27650 206100 27850
rect 205900 27620 206100 27650
rect 206400 27850 206600 27880
rect 206400 27650 206410 27850
rect 206480 27650 206520 27850
rect 206590 27650 206600 27850
rect 206400 27620 206600 27650
rect 206900 27850 207100 27880
rect 206900 27650 206910 27850
rect 206980 27650 207020 27850
rect 207090 27650 207100 27850
rect 206900 27620 207100 27650
rect 207400 27850 207600 27880
rect 207400 27650 207410 27850
rect 207480 27650 207520 27850
rect 207590 27650 207600 27850
rect 207400 27620 207600 27650
rect 207900 27850 208000 27880
rect 207900 27650 207910 27850
rect 207980 27650 208000 27850
rect 207900 27620 208000 27650
rect 204000 27600 204120 27620
rect 204380 27600 204620 27620
rect 204880 27600 205120 27620
rect 205380 27600 205620 27620
rect 205880 27600 206120 27620
rect 206380 27600 206620 27620
rect 206880 27600 207120 27620
rect 207380 27600 207620 27620
rect 207880 27600 208000 27620
rect 204000 27590 208000 27600
rect 204000 27520 204150 27590
rect 204350 27520 204650 27590
rect 204850 27520 205150 27590
rect 205350 27520 205650 27590
rect 205850 27520 206150 27590
rect 206350 27520 206650 27590
rect 206850 27520 207150 27590
rect 207350 27520 207650 27590
rect 207850 27520 208000 27590
rect 204000 27480 208000 27520
rect 204000 27410 204150 27480
rect 204350 27410 204650 27480
rect 204850 27410 205150 27480
rect 205350 27410 205650 27480
rect 205850 27410 206150 27480
rect 206350 27410 206650 27480
rect 206850 27410 207150 27480
rect 207350 27410 207650 27480
rect 207850 27410 208000 27480
rect 204000 27400 208000 27410
rect 204000 27380 204120 27400
rect 204380 27380 204620 27400
rect 204880 27380 205120 27400
rect 205380 27380 205620 27400
rect 205880 27380 206120 27400
rect 206380 27380 206620 27400
rect 206880 27380 207120 27400
rect 207380 27380 207620 27400
rect 207880 27380 208000 27400
rect 204000 27350 204100 27380
rect 204000 27150 204020 27350
rect 204090 27150 204100 27350
rect 204000 27120 204100 27150
rect 204400 27350 204600 27380
rect 204400 27150 204410 27350
rect 204480 27150 204520 27350
rect 204590 27150 204600 27350
rect 204400 27120 204600 27150
rect 204900 27350 205100 27380
rect 204900 27150 204910 27350
rect 204980 27150 205020 27350
rect 205090 27150 205100 27350
rect 204900 27120 205100 27150
rect 205400 27350 205600 27380
rect 205400 27150 205410 27350
rect 205480 27150 205520 27350
rect 205590 27150 205600 27350
rect 205400 27120 205600 27150
rect 205900 27350 206100 27380
rect 205900 27150 205910 27350
rect 205980 27150 206020 27350
rect 206090 27150 206100 27350
rect 205900 27120 206100 27150
rect 206400 27350 206600 27380
rect 206400 27150 206410 27350
rect 206480 27150 206520 27350
rect 206590 27150 206600 27350
rect 206400 27120 206600 27150
rect 206900 27350 207100 27380
rect 206900 27150 206910 27350
rect 206980 27150 207020 27350
rect 207090 27150 207100 27350
rect 206900 27120 207100 27150
rect 207400 27350 207600 27380
rect 207400 27150 207410 27350
rect 207480 27150 207520 27350
rect 207590 27150 207600 27350
rect 207400 27120 207600 27150
rect 207900 27350 208000 27380
rect 207900 27150 207910 27350
rect 207980 27150 208000 27350
rect 207900 27120 208000 27150
rect 204000 27100 204120 27120
rect 204380 27100 204620 27120
rect 204880 27100 205120 27120
rect 205380 27100 205620 27120
rect 205880 27100 206120 27120
rect 206380 27100 206620 27120
rect 206880 27100 207120 27120
rect 207380 27100 207620 27120
rect 207880 27100 208000 27120
rect 204000 27090 208000 27100
rect 204000 27020 204150 27090
rect 204350 27020 204650 27090
rect 204850 27020 205150 27090
rect 205350 27020 205650 27090
rect 205850 27020 206150 27090
rect 206350 27020 206650 27090
rect 206850 27020 207150 27090
rect 207350 27020 207650 27090
rect 207850 27020 208000 27090
rect 204000 26980 208000 27020
rect 204000 26910 204150 26980
rect 204350 26910 204650 26980
rect 204850 26910 205150 26980
rect 205350 26910 205650 26980
rect 205850 26910 206150 26980
rect 206350 26910 206650 26980
rect 206850 26910 207150 26980
rect 207350 26910 207650 26980
rect 207850 26910 208000 26980
rect 204000 26900 208000 26910
rect 204000 26880 204120 26900
rect 204380 26880 204620 26900
rect 204880 26880 205120 26900
rect 205380 26880 205620 26900
rect 205880 26880 206120 26900
rect 206380 26880 206620 26900
rect 206880 26880 207120 26900
rect 207380 26880 207620 26900
rect 207880 26880 208000 26900
rect 204000 26850 204100 26880
rect 204000 26650 204020 26850
rect 204090 26650 204100 26850
rect 204000 26620 204100 26650
rect 204400 26850 204600 26880
rect 204400 26650 204410 26850
rect 204480 26650 204520 26850
rect 204590 26650 204600 26850
rect 204400 26620 204600 26650
rect 204900 26850 205100 26880
rect 204900 26650 204910 26850
rect 204980 26650 205020 26850
rect 205090 26650 205100 26850
rect 204900 26620 205100 26650
rect 205400 26850 205600 26880
rect 205400 26650 205410 26850
rect 205480 26650 205520 26850
rect 205590 26650 205600 26850
rect 205400 26620 205600 26650
rect 205900 26850 206100 26880
rect 205900 26650 205910 26850
rect 205980 26650 206020 26850
rect 206090 26650 206100 26850
rect 205900 26620 206100 26650
rect 206400 26850 206600 26880
rect 206400 26650 206410 26850
rect 206480 26650 206520 26850
rect 206590 26650 206600 26850
rect 206400 26620 206600 26650
rect 206900 26850 207100 26880
rect 206900 26650 206910 26850
rect 206980 26650 207020 26850
rect 207090 26650 207100 26850
rect 206900 26620 207100 26650
rect 207400 26850 207600 26880
rect 207400 26650 207410 26850
rect 207480 26650 207520 26850
rect 207590 26650 207600 26850
rect 207400 26620 207600 26650
rect 207900 26850 208000 26880
rect 207900 26650 207910 26850
rect 207980 26650 208000 26850
rect 207900 26620 208000 26650
rect 204000 26600 204120 26620
rect 204380 26600 204620 26620
rect 204880 26600 205120 26620
rect 205380 26600 205620 26620
rect 205880 26600 206120 26620
rect 206380 26600 206620 26620
rect 206880 26600 207120 26620
rect 207380 26600 207620 26620
rect 207880 26600 208000 26620
rect 204000 26590 208000 26600
rect 204000 26520 204150 26590
rect 204350 26520 204650 26590
rect 204850 26520 205150 26590
rect 205350 26520 205650 26590
rect 205850 26520 206150 26590
rect 206350 26520 206650 26590
rect 206850 26520 207150 26590
rect 207350 26520 207650 26590
rect 207850 26520 208000 26590
rect 204000 26480 208000 26520
rect 204000 26410 204150 26480
rect 204350 26410 204650 26480
rect 204850 26410 205150 26480
rect 205350 26410 205650 26480
rect 205850 26410 206150 26480
rect 206350 26410 206650 26480
rect 206850 26410 207150 26480
rect 207350 26410 207650 26480
rect 207850 26410 208000 26480
rect 204000 26400 208000 26410
rect 204000 26380 204120 26400
rect 204380 26380 204620 26400
rect 204880 26380 205120 26400
rect 205380 26380 205620 26400
rect 205880 26380 206120 26400
rect 206380 26380 206620 26400
rect 206880 26380 207120 26400
rect 207380 26380 207620 26400
rect 207880 26380 208000 26400
rect 204000 26350 204100 26380
rect 204000 26150 204020 26350
rect 204090 26150 204100 26350
rect 204000 26120 204100 26150
rect 204400 26350 204600 26380
rect 204400 26150 204410 26350
rect 204480 26150 204520 26350
rect 204590 26150 204600 26350
rect 204400 26120 204600 26150
rect 204900 26350 205100 26380
rect 204900 26150 204910 26350
rect 204980 26150 205020 26350
rect 205090 26150 205100 26350
rect 204900 26120 205100 26150
rect 205400 26350 205600 26380
rect 205400 26150 205410 26350
rect 205480 26150 205520 26350
rect 205590 26150 205600 26350
rect 205400 26120 205600 26150
rect 205900 26350 206100 26380
rect 205900 26150 205910 26350
rect 205980 26150 206020 26350
rect 206090 26150 206100 26350
rect 205900 26120 206100 26150
rect 206400 26350 206600 26380
rect 206400 26150 206410 26350
rect 206480 26150 206520 26350
rect 206590 26150 206600 26350
rect 206400 26120 206600 26150
rect 206900 26350 207100 26380
rect 206900 26150 206910 26350
rect 206980 26150 207020 26350
rect 207090 26150 207100 26350
rect 206900 26120 207100 26150
rect 207400 26350 207600 26380
rect 207400 26150 207410 26350
rect 207480 26150 207520 26350
rect 207590 26150 207600 26350
rect 207400 26120 207600 26150
rect 207900 26350 208000 26380
rect 207900 26150 207910 26350
rect 207980 26150 208000 26350
rect 207900 26120 208000 26150
rect 204000 26100 204120 26120
rect 204380 26100 204620 26120
rect 204880 26100 205120 26120
rect 205380 26100 205620 26120
rect 205880 26100 206120 26120
rect 206380 26100 206620 26120
rect 206880 26100 207120 26120
rect 207380 26100 207620 26120
rect 207880 26100 208000 26120
rect 204000 26090 208000 26100
rect 204000 26020 204150 26090
rect 204350 26020 204650 26090
rect 204850 26020 205150 26090
rect 205350 26020 205650 26090
rect 205850 26020 206150 26090
rect 206350 26020 206650 26090
rect 206850 26020 207150 26090
rect 207350 26020 207650 26090
rect 207850 26020 208000 26090
rect 204000 25980 208000 26020
rect 204000 25910 204150 25980
rect 204350 25910 204650 25980
rect 204850 25910 205150 25980
rect 205350 25910 205650 25980
rect 205850 25910 206150 25980
rect 206350 25910 206650 25980
rect 206850 25910 207150 25980
rect 207350 25910 207650 25980
rect 207850 25910 208000 25980
rect 204000 25900 208000 25910
rect 204000 25880 204120 25900
rect 204380 25880 204620 25900
rect 204880 25880 205120 25900
rect 205380 25880 205620 25900
rect 205880 25880 206120 25900
rect 206380 25880 206620 25900
rect 206880 25880 207120 25900
rect 207380 25880 207620 25900
rect 207880 25880 208000 25900
rect 204000 25850 204100 25880
rect 204000 25650 204020 25850
rect 204090 25650 204100 25850
rect 204000 25620 204100 25650
rect 204400 25850 204600 25880
rect 204400 25650 204410 25850
rect 204480 25650 204520 25850
rect 204590 25650 204600 25850
rect 204400 25620 204600 25650
rect 204900 25850 205100 25880
rect 204900 25650 204910 25850
rect 204980 25650 205020 25850
rect 205090 25650 205100 25850
rect 204900 25620 205100 25650
rect 205400 25850 205600 25880
rect 205400 25650 205410 25850
rect 205480 25650 205520 25850
rect 205590 25650 205600 25850
rect 205400 25620 205600 25650
rect 205900 25850 206100 25880
rect 205900 25650 205910 25850
rect 205980 25650 206020 25850
rect 206090 25650 206100 25850
rect 205900 25620 206100 25650
rect 206400 25850 206600 25880
rect 206400 25650 206410 25850
rect 206480 25650 206520 25850
rect 206590 25650 206600 25850
rect 206400 25620 206600 25650
rect 206900 25850 207100 25880
rect 206900 25650 206910 25850
rect 206980 25650 207020 25850
rect 207090 25650 207100 25850
rect 206900 25620 207100 25650
rect 207400 25850 207600 25880
rect 207400 25650 207410 25850
rect 207480 25650 207520 25850
rect 207590 25650 207600 25850
rect 207400 25620 207600 25650
rect 207900 25850 208000 25880
rect 207900 25650 207910 25850
rect 207980 25650 208000 25850
rect 207900 25620 208000 25650
rect 204000 25600 204120 25620
rect 204380 25600 204620 25620
rect 204880 25600 205120 25620
rect 205380 25600 205620 25620
rect 205880 25600 206120 25620
rect 206380 25600 206620 25620
rect 206880 25600 207120 25620
rect 207380 25600 207620 25620
rect 207880 25600 208000 25620
rect 204000 25590 208000 25600
rect 204000 25520 204150 25590
rect 204350 25520 204650 25590
rect 204850 25520 205150 25590
rect 205350 25520 205650 25590
rect 205850 25520 206150 25590
rect 206350 25520 206650 25590
rect 206850 25520 207150 25590
rect 207350 25520 207650 25590
rect 207850 25520 208000 25590
rect 204000 25480 208000 25520
rect 204000 25410 204150 25480
rect 204350 25410 204650 25480
rect 204850 25410 205150 25480
rect 205350 25410 205650 25480
rect 205850 25410 206150 25480
rect 206350 25410 206650 25480
rect 206850 25410 207150 25480
rect 207350 25410 207650 25480
rect 207850 25410 208000 25480
rect 204000 25400 208000 25410
rect 204000 25380 204120 25400
rect 204380 25380 204620 25400
rect 204880 25380 205120 25400
rect 205380 25380 205620 25400
rect 205880 25380 206120 25400
rect 206380 25380 206620 25400
rect 206880 25380 207120 25400
rect 207380 25380 207620 25400
rect 207880 25380 208000 25400
rect 204000 25350 204100 25380
rect 204000 25150 204020 25350
rect 204090 25150 204100 25350
rect 204000 25120 204100 25150
rect 204400 25350 204600 25380
rect 204400 25150 204410 25350
rect 204480 25150 204520 25350
rect 204590 25150 204600 25350
rect 204400 25120 204600 25150
rect 204900 25350 205100 25380
rect 204900 25150 204910 25350
rect 204980 25150 205020 25350
rect 205090 25150 205100 25350
rect 204900 25120 205100 25150
rect 205400 25350 205600 25380
rect 205400 25150 205410 25350
rect 205480 25150 205520 25350
rect 205590 25150 205600 25350
rect 205400 25120 205600 25150
rect 205900 25350 206100 25380
rect 205900 25150 205910 25350
rect 205980 25150 206020 25350
rect 206090 25150 206100 25350
rect 205900 25120 206100 25150
rect 206400 25350 206600 25380
rect 206400 25150 206410 25350
rect 206480 25150 206520 25350
rect 206590 25150 206600 25350
rect 206400 25120 206600 25150
rect 206900 25350 207100 25380
rect 206900 25150 206910 25350
rect 206980 25150 207020 25350
rect 207090 25150 207100 25350
rect 206900 25120 207100 25150
rect 207400 25350 207600 25380
rect 207400 25150 207410 25350
rect 207480 25150 207520 25350
rect 207590 25150 207600 25350
rect 207400 25120 207600 25150
rect 207900 25350 208000 25380
rect 207900 25150 207910 25350
rect 207980 25150 208000 25350
rect 207900 25120 208000 25150
rect 204000 25100 204120 25120
rect 204380 25100 204620 25120
rect 204880 25100 205120 25120
rect 205380 25100 205620 25120
rect 205880 25100 206120 25120
rect 206380 25100 206620 25120
rect 206880 25100 207120 25120
rect 207380 25100 207620 25120
rect 207880 25100 208000 25120
rect 204000 25090 208000 25100
rect 204000 25020 204150 25090
rect 204350 25020 204650 25090
rect 204850 25020 205150 25090
rect 205350 25020 205650 25090
rect 205850 25020 206150 25090
rect 206350 25020 206650 25090
rect 206850 25020 207150 25090
rect 207350 25020 207650 25090
rect 207850 25020 208000 25090
rect 204000 24980 208000 25020
rect 204000 24910 204150 24980
rect 204350 24910 204650 24980
rect 204850 24910 205150 24980
rect 205350 24910 205650 24980
rect 205850 24910 206150 24980
rect 206350 24910 206650 24980
rect 206850 24910 207150 24980
rect 207350 24910 207650 24980
rect 207850 24910 208000 24980
rect 204000 24900 208000 24910
rect 204000 24880 204120 24900
rect 204380 24880 204620 24900
rect 204880 24880 205120 24900
rect 205380 24880 205620 24900
rect 205880 24880 206120 24900
rect 206380 24880 206620 24900
rect 206880 24880 207120 24900
rect 207380 24880 207620 24900
rect 207880 24880 208000 24900
rect 204000 24850 204100 24880
rect 204000 24650 204020 24850
rect 204090 24650 204100 24850
rect 204000 24620 204100 24650
rect 204400 24850 204600 24880
rect 204400 24650 204410 24850
rect 204480 24650 204520 24850
rect 204590 24650 204600 24850
rect 204400 24620 204600 24650
rect 204900 24850 205100 24880
rect 204900 24650 204910 24850
rect 204980 24650 205020 24850
rect 205090 24650 205100 24850
rect 204900 24620 205100 24650
rect 205400 24850 205600 24880
rect 205400 24650 205410 24850
rect 205480 24650 205520 24850
rect 205590 24650 205600 24850
rect 205400 24620 205600 24650
rect 205900 24850 206100 24880
rect 205900 24650 205910 24850
rect 205980 24650 206020 24850
rect 206090 24650 206100 24850
rect 205900 24620 206100 24650
rect 206400 24850 206600 24880
rect 206400 24650 206410 24850
rect 206480 24650 206520 24850
rect 206590 24650 206600 24850
rect 206400 24620 206600 24650
rect 206900 24850 207100 24880
rect 206900 24650 206910 24850
rect 206980 24650 207020 24850
rect 207090 24650 207100 24850
rect 206900 24620 207100 24650
rect 207400 24850 207600 24880
rect 207400 24650 207410 24850
rect 207480 24650 207520 24850
rect 207590 24650 207600 24850
rect 207400 24620 207600 24650
rect 207900 24850 208000 24880
rect 207900 24650 207910 24850
rect 207980 24650 208000 24850
rect 207900 24620 208000 24650
rect 204000 24600 204120 24620
rect 204380 24600 204620 24620
rect 204880 24600 205120 24620
rect 205380 24600 205620 24620
rect 205880 24600 206120 24620
rect 206380 24600 206620 24620
rect 206880 24600 207120 24620
rect 207380 24600 207620 24620
rect 207880 24600 208000 24620
rect 204000 24590 208000 24600
rect 204000 24520 204150 24590
rect 204350 24520 204650 24590
rect 204850 24520 205150 24590
rect 205350 24520 205650 24590
rect 205850 24520 206150 24590
rect 206350 24520 206650 24590
rect 206850 24520 207150 24590
rect 207350 24520 207650 24590
rect 207850 24520 208000 24590
rect 204000 24480 208000 24520
rect 204000 24410 204150 24480
rect 204350 24410 204650 24480
rect 204850 24410 205150 24480
rect 205350 24410 205650 24480
rect 205850 24410 206150 24480
rect 206350 24410 206650 24480
rect 206850 24410 207150 24480
rect 207350 24410 207650 24480
rect 207850 24410 208000 24480
rect 204000 24400 208000 24410
rect 204000 24380 204120 24400
rect 204380 24380 204620 24400
rect 204880 24380 205120 24400
rect 205380 24380 205620 24400
rect 205880 24380 206120 24400
rect 206380 24380 206620 24400
rect 206880 24380 207120 24400
rect 207380 24380 207620 24400
rect 207880 24380 208000 24400
rect 204000 24350 204100 24380
rect 204000 24150 204020 24350
rect 204090 24150 204100 24350
rect 204000 24120 204100 24150
rect 204400 24350 204600 24380
rect 204400 24150 204410 24350
rect 204480 24150 204520 24350
rect 204590 24150 204600 24350
rect 204400 24120 204600 24150
rect 204900 24350 205100 24380
rect 204900 24150 204910 24350
rect 204980 24150 205020 24350
rect 205090 24150 205100 24350
rect 204900 24120 205100 24150
rect 205400 24350 205600 24380
rect 205400 24150 205410 24350
rect 205480 24150 205520 24350
rect 205590 24150 205600 24350
rect 205400 24120 205600 24150
rect 205900 24350 206100 24380
rect 205900 24150 205910 24350
rect 205980 24150 206020 24350
rect 206090 24150 206100 24350
rect 205900 24120 206100 24150
rect 206400 24350 206600 24380
rect 206400 24150 206410 24350
rect 206480 24150 206520 24350
rect 206590 24150 206600 24350
rect 206400 24120 206600 24150
rect 206900 24350 207100 24380
rect 206900 24150 206910 24350
rect 206980 24150 207020 24350
rect 207090 24150 207100 24350
rect 206900 24120 207100 24150
rect 207400 24350 207600 24380
rect 207400 24150 207410 24350
rect 207480 24150 207520 24350
rect 207590 24150 207600 24350
rect 207400 24120 207600 24150
rect 207900 24350 208000 24380
rect 207900 24150 207910 24350
rect 207980 24150 208000 24350
rect 207900 24120 208000 24150
rect 204000 24100 204120 24120
rect 204380 24100 204620 24120
rect 204880 24100 205120 24120
rect 205380 24100 205620 24120
rect 205880 24100 206120 24120
rect 206380 24100 206620 24120
rect 206880 24100 207120 24120
rect 207380 24100 207620 24120
rect 207880 24100 208000 24120
rect 204000 24090 208000 24100
rect 204000 24020 204150 24090
rect 204350 24020 204650 24090
rect 204850 24020 205150 24090
rect 205350 24020 205650 24090
rect 205850 24020 206150 24090
rect 206350 24020 206650 24090
rect 206850 24020 207150 24090
rect 207350 24020 207650 24090
rect 207850 24020 208000 24090
rect 204000 23980 208000 24020
rect 204000 23910 204150 23980
rect 204350 23910 204650 23980
rect 204850 23910 205150 23980
rect 205350 23910 205650 23980
rect 205850 23910 206150 23980
rect 206350 23910 206650 23980
rect 206850 23910 207150 23980
rect 207350 23910 207650 23980
rect 207850 23910 208000 23980
rect 204000 23900 208000 23910
rect 204000 23880 204120 23900
rect 204380 23880 204620 23900
rect 204880 23880 205120 23900
rect 205380 23880 205620 23900
rect 205880 23880 206120 23900
rect 206380 23880 206620 23900
rect 206880 23880 207120 23900
rect 207380 23880 207620 23900
rect 207880 23880 208000 23900
rect 204000 23850 204100 23880
rect 204000 23650 204020 23850
rect 204090 23650 204100 23850
rect 204000 23620 204100 23650
rect 204400 23850 204600 23880
rect 204400 23650 204410 23850
rect 204480 23650 204520 23850
rect 204590 23650 204600 23850
rect 204400 23620 204600 23650
rect 204900 23850 205100 23880
rect 204900 23650 204910 23850
rect 204980 23650 205020 23850
rect 205090 23650 205100 23850
rect 204900 23620 205100 23650
rect 205400 23850 205600 23880
rect 205400 23650 205410 23850
rect 205480 23650 205520 23850
rect 205590 23650 205600 23850
rect 205400 23620 205600 23650
rect 205900 23850 206100 23880
rect 205900 23650 205910 23850
rect 205980 23650 206020 23850
rect 206090 23650 206100 23850
rect 205900 23620 206100 23650
rect 206400 23850 206600 23880
rect 206400 23650 206410 23850
rect 206480 23650 206520 23850
rect 206590 23650 206600 23850
rect 206400 23620 206600 23650
rect 206900 23850 207100 23880
rect 206900 23650 206910 23850
rect 206980 23650 207020 23850
rect 207090 23650 207100 23850
rect 206900 23620 207100 23650
rect 207400 23850 207600 23880
rect 207400 23650 207410 23850
rect 207480 23650 207520 23850
rect 207590 23650 207600 23850
rect 207400 23620 207600 23650
rect 207900 23850 208000 23880
rect 207900 23650 207910 23850
rect 207980 23650 208000 23850
rect 207900 23620 208000 23650
rect 204000 23600 204120 23620
rect 204380 23600 204620 23620
rect 204880 23600 205120 23620
rect 205380 23600 205620 23620
rect 205880 23600 206120 23620
rect 206380 23600 206620 23620
rect 206880 23600 207120 23620
rect 207380 23600 207620 23620
rect 207880 23600 208000 23620
rect 204000 23590 208000 23600
rect 204000 23520 204150 23590
rect 204350 23520 204650 23590
rect 204850 23520 205150 23590
rect 205350 23520 205650 23590
rect 205850 23520 206150 23590
rect 206350 23520 206650 23590
rect 206850 23520 207150 23590
rect 207350 23520 207650 23590
rect 207850 23520 208000 23590
rect 204000 23480 208000 23520
rect 204000 23410 204150 23480
rect 204350 23410 204650 23480
rect 204850 23410 205150 23480
rect 205350 23410 205650 23480
rect 205850 23410 206150 23480
rect 206350 23410 206650 23480
rect 206850 23410 207150 23480
rect 207350 23410 207650 23480
rect 207850 23410 208000 23480
rect 204000 23400 208000 23410
rect 204000 23380 204120 23400
rect 204380 23380 204620 23400
rect 204880 23380 205120 23400
rect 205380 23380 205620 23400
rect 205880 23380 206120 23400
rect 206380 23380 206620 23400
rect 206880 23380 207120 23400
rect 207380 23380 207620 23400
rect 207880 23380 208000 23400
rect 204000 23350 204100 23380
rect 204000 23150 204020 23350
rect 204090 23150 204100 23350
rect 204000 23120 204100 23150
rect 204400 23350 204600 23380
rect 204400 23150 204410 23350
rect 204480 23150 204520 23350
rect 204590 23150 204600 23350
rect 204400 23120 204600 23150
rect 204900 23350 205100 23380
rect 204900 23150 204910 23350
rect 204980 23150 205020 23350
rect 205090 23150 205100 23350
rect 204900 23120 205100 23150
rect 205400 23350 205600 23380
rect 205400 23150 205410 23350
rect 205480 23150 205520 23350
rect 205590 23150 205600 23350
rect 205400 23120 205600 23150
rect 205900 23350 206100 23380
rect 205900 23150 205910 23350
rect 205980 23150 206020 23350
rect 206090 23150 206100 23350
rect 205900 23120 206100 23150
rect 206400 23350 206600 23380
rect 206400 23150 206410 23350
rect 206480 23150 206520 23350
rect 206590 23150 206600 23350
rect 206400 23120 206600 23150
rect 206900 23350 207100 23380
rect 206900 23150 206910 23350
rect 206980 23150 207020 23350
rect 207090 23150 207100 23350
rect 206900 23120 207100 23150
rect 207400 23350 207600 23380
rect 207400 23150 207410 23350
rect 207480 23150 207520 23350
rect 207590 23150 207600 23350
rect 207400 23120 207600 23150
rect 207900 23350 208000 23380
rect 207900 23150 207910 23350
rect 207980 23150 208000 23350
rect 207900 23120 208000 23150
rect 204000 23100 204120 23120
rect 204380 23100 204620 23120
rect 204880 23100 205120 23120
rect 205380 23100 205620 23120
rect 205880 23100 206120 23120
rect 206380 23100 206620 23120
rect 206880 23100 207120 23120
rect 207380 23100 207620 23120
rect 207880 23100 208000 23120
rect 204000 23090 208000 23100
rect 204000 23020 204150 23090
rect 204350 23020 204650 23090
rect 204850 23020 205150 23090
rect 205350 23020 205650 23090
rect 205850 23020 206150 23090
rect 206350 23020 206650 23090
rect 206850 23020 207150 23090
rect 207350 23020 207650 23090
rect 207850 23020 208000 23090
rect 204000 22980 208000 23020
rect 204000 22910 204150 22980
rect 204350 22910 204650 22980
rect 204850 22910 205150 22980
rect 205350 22910 205650 22980
rect 205850 22910 206150 22980
rect 206350 22910 206650 22980
rect 206850 22910 207150 22980
rect 207350 22910 207650 22980
rect 207850 22910 208000 22980
rect 204000 22900 208000 22910
rect 204000 22880 204120 22900
rect 204380 22880 204620 22900
rect 204880 22880 205120 22900
rect 205380 22880 205620 22900
rect 205880 22880 206120 22900
rect 206380 22880 206620 22900
rect 206880 22880 207120 22900
rect 207380 22880 207620 22900
rect 207880 22880 208000 22900
rect 204000 22850 204100 22880
rect 204000 22650 204020 22850
rect 204090 22650 204100 22850
rect 204000 22620 204100 22650
rect 204400 22850 204600 22880
rect 204400 22650 204410 22850
rect 204480 22650 204520 22850
rect 204590 22650 204600 22850
rect 204400 22620 204600 22650
rect 204900 22850 205100 22880
rect 204900 22650 204910 22850
rect 204980 22650 205020 22850
rect 205090 22650 205100 22850
rect 204900 22620 205100 22650
rect 205400 22850 205600 22880
rect 205400 22650 205410 22850
rect 205480 22650 205520 22850
rect 205590 22650 205600 22850
rect 205400 22620 205600 22650
rect 205900 22850 206100 22880
rect 205900 22650 205910 22850
rect 205980 22650 206020 22850
rect 206090 22650 206100 22850
rect 205900 22620 206100 22650
rect 206400 22850 206600 22880
rect 206400 22650 206410 22850
rect 206480 22650 206520 22850
rect 206590 22650 206600 22850
rect 206400 22620 206600 22650
rect 206900 22850 207100 22880
rect 206900 22650 206910 22850
rect 206980 22650 207020 22850
rect 207090 22650 207100 22850
rect 206900 22620 207100 22650
rect 207400 22850 207600 22880
rect 207400 22650 207410 22850
rect 207480 22650 207520 22850
rect 207590 22650 207600 22850
rect 207400 22620 207600 22650
rect 207900 22850 208000 22880
rect 207900 22650 207910 22850
rect 207980 22650 208000 22850
rect 207900 22620 208000 22650
rect 204000 22600 204120 22620
rect 204380 22600 204620 22620
rect 204880 22600 205120 22620
rect 205380 22600 205620 22620
rect 205880 22600 206120 22620
rect 206380 22600 206620 22620
rect 206880 22600 207120 22620
rect 207380 22600 207620 22620
rect 207880 22600 208000 22620
rect 204000 22590 208000 22600
rect 204000 22520 204150 22590
rect 204350 22520 204650 22590
rect 204850 22520 205150 22590
rect 205350 22520 205650 22590
rect 205850 22520 206150 22590
rect 206350 22520 206650 22590
rect 206850 22520 207150 22590
rect 207350 22520 207650 22590
rect 207850 22520 208000 22590
rect 204000 22480 208000 22520
rect 204000 22410 204150 22480
rect 204350 22410 204650 22480
rect 204850 22410 205150 22480
rect 205350 22410 205650 22480
rect 205850 22410 206150 22480
rect 206350 22410 206650 22480
rect 206850 22410 207150 22480
rect 207350 22410 207650 22480
rect 207850 22410 208000 22480
rect 204000 22400 208000 22410
rect 204000 22380 204120 22400
rect 204380 22380 204620 22400
rect 204880 22380 205120 22400
rect 205380 22380 205620 22400
rect 205880 22380 206120 22400
rect 206380 22380 206620 22400
rect 206880 22380 207120 22400
rect 207380 22380 207620 22400
rect 207880 22380 208000 22400
rect 204000 22350 204100 22380
rect 204000 22150 204020 22350
rect 204090 22150 204100 22350
rect 204000 22120 204100 22150
rect 204400 22350 204600 22380
rect 204400 22150 204410 22350
rect 204480 22150 204520 22350
rect 204590 22150 204600 22350
rect 204400 22120 204600 22150
rect 204900 22350 205100 22380
rect 204900 22150 204910 22350
rect 204980 22150 205020 22350
rect 205090 22150 205100 22350
rect 204900 22120 205100 22150
rect 205400 22350 205600 22380
rect 205400 22150 205410 22350
rect 205480 22150 205520 22350
rect 205590 22150 205600 22350
rect 205400 22120 205600 22150
rect 205900 22350 206100 22380
rect 205900 22150 205910 22350
rect 205980 22150 206020 22350
rect 206090 22150 206100 22350
rect 205900 22120 206100 22150
rect 206400 22350 206600 22380
rect 206400 22150 206410 22350
rect 206480 22150 206520 22350
rect 206590 22150 206600 22350
rect 206400 22120 206600 22150
rect 206900 22350 207100 22380
rect 206900 22150 206910 22350
rect 206980 22150 207020 22350
rect 207090 22150 207100 22350
rect 206900 22120 207100 22150
rect 207400 22350 207600 22380
rect 207400 22150 207410 22350
rect 207480 22150 207520 22350
rect 207590 22150 207600 22350
rect 207400 22120 207600 22150
rect 207900 22350 208000 22380
rect 207900 22150 207910 22350
rect 207980 22150 208000 22350
rect 207900 22120 208000 22150
rect 204000 22100 204120 22120
rect 204380 22100 204620 22120
rect 204880 22100 205120 22120
rect 205380 22100 205620 22120
rect 205880 22100 206120 22120
rect 206380 22100 206620 22120
rect 206880 22100 207120 22120
rect 207380 22100 207620 22120
rect 207880 22100 208000 22120
rect 204000 22090 208000 22100
rect 204000 22020 204150 22090
rect 204350 22020 204650 22090
rect 204850 22020 205150 22090
rect 205350 22020 205650 22090
rect 205850 22020 206150 22090
rect 206350 22020 206650 22090
rect 206850 22020 207150 22090
rect 207350 22020 207650 22090
rect 207850 22020 208000 22090
rect 204000 21980 208000 22020
rect 204000 21910 204150 21980
rect 204350 21910 204650 21980
rect 204850 21910 205150 21980
rect 205350 21910 205650 21980
rect 205850 21910 206150 21980
rect 206350 21910 206650 21980
rect 206850 21910 207150 21980
rect 207350 21910 207650 21980
rect 207850 21910 208000 21980
rect 204000 21900 208000 21910
rect 204000 21880 204120 21900
rect 204380 21880 204620 21900
rect 204880 21880 205120 21900
rect 205380 21880 205620 21900
rect 205880 21880 206120 21900
rect 206380 21880 206620 21900
rect 206880 21880 207120 21900
rect 207380 21880 207620 21900
rect 207880 21880 208000 21900
rect 204000 21850 204100 21880
rect 204000 21650 204020 21850
rect 204090 21650 204100 21850
rect 204000 21620 204100 21650
rect 204400 21850 204600 21880
rect 204400 21650 204410 21850
rect 204480 21650 204520 21850
rect 204590 21650 204600 21850
rect 204400 21620 204600 21650
rect 204900 21850 205100 21880
rect 204900 21650 204910 21850
rect 204980 21650 205020 21850
rect 205090 21650 205100 21850
rect 204900 21620 205100 21650
rect 205400 21850 205600 21880
rect 205400 21650 205410 21850
rect 205480 21650 205520 21850
rect 205590 21650 205600 21850
rect 205400 21620 205600 21650
rect 205900 21850 206100 21880
rect 205900 21650 205910 21850
rect 205980 21650 206020 21850
rect 206090 21650 206100 21850
rect 205900 21620 206100 21650
rect 206400 21850 206600 21880
rect 206400 21650 206410 21850
rect 206480 21650 206520 21850
rect 206590 21650 206600 21850
rect 206400 21620 206600 21650
rect 206900 21850 207100 21880
rect 206900 21650 206910 21850
rect 206980 21650 207020 21850
rect 207090 21650 207100 21850
rect 206900 21620 207100 21650
rect 207400 21850 207600 21880
rect 207400 21650 207410 21850
rect 207480 21650 207520 21850
rect 207590 21650 207600 21850
rect 207400 21620 207600 21650
rect 207900 21850 208000 21880
rect 207900 21650 207910 21850
rect 207980 21650 208000 21850
rect 207900 21620 208000 21650
rect 204000 21600 204120 21620
rect 204380 21600 204620 21620
rect 204880 21600 205120 21620
rect 205380 21600 205620 21620
rect 205880 21600 206120 21620
rect 206380 21600 206620 21620
rect 206880 21600 207120 21620
rect 207380 21600 207620 21620
rect 207880 21600 208000 21620
rect 204000 21590 208000 21600
rect 204000 21520 204150 21590
rect 204350 21520 204650 21590
rect 204850 21520 205150 21590
rect 205350 21520 205650 21590
rect 205850 21520 206150 21590
rect 206350 21520 206650 21590
rect 206850 21520 207150 21590
rect 207350 21520 207650 21590
rect 207850 21520 208000 21590
rect 204000 21480 208000 21520
rect 204000 21410 204150 21480
rect 204350 21410 204650 21480
rect 204850 21410 205150 21480
rect 205350 21410 205650 21480
rect 205850 21410 206150 21480
rect 206350 21410 206650 21480
rect 206850 21410 207150 21480
rect 207350 21410 207650 21480
rect 207850 21410 208000 21480
rect 204000 21400 208000 21410
rect 204000 21380 204120 21400
rect 204380 21380 204620 21400
rect 204880 21380 205120 21400
rect 205380 21380 205620 21400
rect 205880 21380 206120 21400
rect 206380 21380 206620 21400
rect 206880 21380 207120 21400
rect 207380 21380 207620 21400
rect 207880 21380 208000 21400
rect 204000 21350 204100 21380
rect 204000 21150 204020 21350
rect 204090 21150 204100 21350
rect 204000 21120 204100 21150
rect 204400 21350 204600 21380
rect 204400 21150 204410 21350
rect 204480 21150 204520 21350
rect 204590 21150 204600 21350
rect 204400 21120 204600 21150
rect 204900 21350 205100 21380
rect 204900 21150 204910 21350
rect 204980 21150 205020 21350
rect 205090 21150 205100 21350
rect 204900 21120 205100 21150
rect 205400 21350 205600 21380
rect 205400 21150 205410 21350
rect 205480 21150 205520 21350
rect 205590 21150 205600 21350
rect 205400 21120 205600 21150
rect 205900 21350 206100 21380
rect 205900 21150 205910 21350
rect 205980 21150 206020 21350
rect 206090 21150 206100 21350
rect 205900 21120 206100 21150
rect 206400 21350 206600 21380
rect 206400 21150 206410 21350
rect 206480 21150 206520 21350
rect 206590 21150 206600 21350
rect 206400 21120 206600 21150
rect 206900 21350 207100 21380
rect 206900 21150 206910 21350
rect 206980 21150 207020 21350
rect 207090 21150 207100 21350
rect 206900 21120 207100 21150
rect 207400 21350 207600 21380
rect 207400 21150 207410 21350
rect 207480 21150 207520 21350
rect 207590 21150 207600 21350
rect 207400 21120 207600 21150
rect 207900 21350 208000 21380
rect 207900 21150 207910 21350
rect 207980 21150 208000 21350
rect 207900 21120 208000 21150
rect 204000 21100 204120 21120
rect 204380 21100 204620 21120
rect 204880 21100 205120 21120
rect 205380 21100 205620 21120
rect 205880 21100 206120 21120
rect 206380 21100 206620 21120
rect 206880 21100 207120 21120
rect 207380 21100 207620 21120
rect 207880 21100 208000 21120
rect 204000 21090 208000 21100
rect 204000 21020 204150 21090
rect 204350 21020 204650 21090
rect 204850 21020 205150 21090
rect 205350 21020 205650 21090
rect 205850 21020 206150 21090
rect 206350 21020 206650 21090
rect 206850 21020 207150 21090
rect 207350 21020 207650 21090
rect 207850 21020 208000 21090
rect 204000 20980 208000 21020
rect 204000 20910 204150 20980
rect 204350 20910 204650 20980
rect 204850 20910 205150 20980
rect 205350 20910 205650 20980
rect 205850 20910 206150 20980
rect 206350 20910 206650 20980
rect 206850 20910 207150 20980
rect 207350 20910 207650 20980
rect 207850 20910 208000 20980
rect 204000 20900 208000 20910
rect 204000 20880 204120 20900
rect 204380 20880 204620 20900
rect 204880 20880 205120 20900
rect 205380 20880 205620 20900
rect 205880 20880 206120 20900
rect 206380 20880 206620 20900
rect 206880 20880 207120 20900
rect 207380 20880 207620 20900
rect 207880 20880 208000 20900
rect 204000 20850 204100 20880
rect 204000 20650 204020 20850
rect 204090 20650 204100 20850
rect 204000 20620 204100 20650
rect 204400 20850 204600 20880
rect 204400 20650 204410 20850
rect 204480 20650 204520 20850
rect 204590 20650 204600 20850
rect 204400 20620 204600 20650
rect 204900 20850 205100 20880
rect 204900 20650 204910 20850
rect 204980 20650 205020 20850
rect 205090 20650 205100 20850
rect 204900 20620 205100 20650
rect 205400 20850 205600 20880
rect 205400 20650 205410 20850
rect 205480 20650 205520 20850
rect 205590 20650 205600 20850
rect 205400 20620 205600 20650
rect 205900 20850 206100 20880
rect 205900 20650 205910 20850
rect 205980 20650 206020 20850
rect 206090 20650 206100 20850
rect 205900 20620 206100 20650
rect 206400 20850 206600 20880
rect 206400 20650 206410 20850
rect 206480 20650 206520 20850
rect 206590 20650 206600 20850
rect 206400 20620 206600 20650
rect 206900 20850 207100 20880
rect 206900 20650 206910 20850
rect 206980 20650 207020 20850
rect 207090 20650 207100 20850
rect 206900 20620 207100 20650
rect 207400 20850 207600 20880
rect 207400 20650 207410 20850
rect 207480 20650 207520 20850
rect 207590 20650 207600 20850
rect 207400 20620 207600 20650
rect 207900 20850 208000 20880
rect 207900 20650 207910 20850
rect 207980 20650 208000 20850
rect 207900 20620 208000 20650
rect 204000 20600 204120 20620
rect 204380 20600 204620 20620
rect 204880 20600 205120 20620
rect 205380 20600 205620 20620
rect 205880 20600 206120 20620
rect 206380 20600 206620 20620
rect 206880 20600 207120 20620
rect 207380 20600 207620 20620
rect 207880 20600 208000 20620
rect 204000 20590 208000 20600
rect 204000 20520 204150 20590
rect 204350 20520 204650 20590
rect 204850 20520 205150 20590
rect 205350 20520 205650 20590
rect 205850 20520 206150 20590
rect 206350 20520 206650 20590
rect 206850 20520 207150 20590
rect 207350 20520 207650 20590
rect 207850 20520 208000 20590
rect 204000 20480 208000 20520
rect 204000 20410 204150 20480
rect 204350 20410 204650 20480
rect 204850 20410 205150 20480
rect 205350 20410 205650 20480
rect 205850 20410 206150 20480
rect 206350 20410 206650 20480
rect 206850 20410 207150 20480
rect 207350 20410 207650 20480
rect 207850 20410 208000 20480
rect 204000 20400 208000 20410
rect 204000 20380 204120 20400
rect 204380 20380 204620 20400
rect 204880 20380 205120 20400
rect 205380 20380 205620 20400
rect 205880 20380 206120 20400
rect 206380 20380 206620 20400
rect 206880 20380 207120 20400
rect 207380 20380 207620 20400
rect 207880 20380 208000 20400
rect 204000 20350 204100 20380
rect 204000 20150 204020 20350
rect 204090 20150 204100 20350
rect 204000 20120 204100 20150
rect 204400 20350 204600 20380
rect 204400 20150 204410 20350
rect 204480 20150 204520 20350
rect 204590 20150 204600 20350
rect 204400 20120 204600 20150
rect 204900 20350 205100 20380
rect 204900 20150 204910 20350
rect 204980 20150 205020 20350
rect 205090 20150 205100 20350
rect 204900 20120 205100 20150
rect 205400 20350 205600 20380
rect 205400 20150 205410 20350
rect 205480 20150 205520 20350
rect 205590 20150 205600 20350
rect 205400 20120 205600 20150
rect 205900 20350 206100 20380
rect 205900 20150 205910 20350
rect 205980 20150 206020 20350
rect 206090 20150 206100 20350
rect 205900 20120 206100 20150
rect 206400 20350 206600 20380
rect 206400 20150 206410 20350
rect 206480 20150 206520 20350
rect 206590 20150 206600 20350
rect 206400 20120 206600 20150
rect 206900 20350 207100 20380
rect 206900 20150 206910 20350
rect 206980 20150 207020 20350
rect 207090 20150 207100 20350
rect 206900 20120 207100 20150
rect 207400 20350 207600 20380
rect 207400 20150 207410 20350
rect 207480 20150 207520 20350
rect 207590 20150 207600 20350
rect 207400 20120 207600 20150
rect 207900 20350 208000 20380
rect 207900 20150 207910 20350
rect 207980 20150 208000 20350
rect 207900 20120 208000 20150
rect 204000 20100 204120 20120
rect 204380 20100 204620 20120
rect 204880 20100 205120 20120
rect 205380 20100 205620 20120
rect 205880 20100 206120 20120
rect 206380 20100 206620 20120
rect 206880 20100 207120 20120
rect 207380 20100 207620 20120
rect 207880 20100 208000 20120
rect 204000 20090 208000 20100
rect 204000 20020 204150 20090
rect 204350 20020 204650 20090
rect 204850 20020 205150 20090
rect 205350 20020 205650 20090
rect 205850 20020 206150 20090
rect 206350 20020 206650 20090
rect 206850 20020 207150 20090
rect 207350 20020 207650 20090
rect 207850 20020 208000 20090
rect 204000 19980 208000 20020
rect 204000 19910 204150 19980
rect 204350 19910 204650 19980
rect 204850 19910 205150 19980
rect 205350 19910 205650 19980
rect 205850 19910 206150 19980
rect 206350 19910 206650 19980
rect 206850 19910 207150 19980
rect 207350 19910 207650 19980
rect 207850 19910 208000 19980
rect 204000 19900 208000 19910
rect 204000 19880 204120 19900
rect 204380 19880 204620 19900
rect 204880 19880 205120 19900
rect 205380 19880 205620 19900
rect 205880 19880 206120 19900
rect 206380 19880 206620 19900
rect 206880 19880 207120 19900
rect 207380 19880 207620 19900
rect 207880 19880 208000 19900
rect 204000 19850 204100 19880
rect 204000 19650 204020 19850
rect 204090 19650 204100 19850
rect 204000 19620 204100 19650
rect 204400 19850 204600 19880
rect 204400 19650 204410 19850
rect 204480 19650 204520 19850
rect 204590 19650 204600 19850
rect 204400 19620 204600 19650
rect 204900 19850 205100 19880
rect 204900 19650 204910 19850
rect 204980 19650 205020 19850
rect 205090 19650 205100 19850
rect 204900 19620 205100 19650
rect 205400 19850 205600 19880
rect 205400 19650 205410 19850
rect 205480 19650 205520 19850
rect 205590 19650 205600 19850
rect 205400 19620 205600 19650
rect 205900 19850 206100 19880
rect 205900 19650 205910 19850
rect 205980 19650 206020 19850
rect 206090 19650 206100 19850
rect 205900 19620 206100 19650
rect 206400 19850 206600 19880
rect 206400 19650 206410 19850
rect 206480 19650 206520 19850
rect 206590 19650 206600 19850
rect 206400 19620 206600 19650
rect 206900 19850 207100 19880
rect 206900 19650 206910 19850
rect 206980 19650 207020 19850
rect 207090 19650 207100 19850
rect 206900 19620 207100 19650
rect 207400 19850 207600 19880
rect 207400 19650 207410 19850
rect 207480 19650 207520 19850
rect 207590 19650 207600 19850
rect 207400 19620 207600 19650
rect 207900 19850 208000 19880
rect 207900 19650 207910 19850
rect 207980 19650 208000 19850
rect 207900 19620 208000 19650
rect 204000 19600 204120 19620
rect 204380 19600 204620 19620
rect 204880 19600 205120 19620
rect 205380 19600 205620 19620
rect 205880 19600 206120 19620
rect 206380 19600 206620 19620
rect 206880 19600 207120 19620
rect 207380 19600 207620 19620
rect 207880 19600 208000 19620
rect 204000 19590 208000 19600
rect 204000 19520 204150 19590
rect 204350 19520 204650 19590
rect 204850 19520 205150 19590
rect 205350 19520 205650 19590
rect 205850 19520 206150 19590
rect 206350 19520 206650 19590
rect 206850 19520 207150 19590
rect 207350 19520 207650 19590
rect 207850 19520 208000 19590
rect 204000 19480 208000 19520
rect 204000 19410 204150 19480
rect 204350 19410 204650 19480
rect 204850 19410 205150 19480
rect 205350 19410 205650 19480
rect 205850 19410 206150 19480
rect 206350 19410 206650 19480
rect 206850 19410 207150 19480
rect 207350 19410 207650 19480
rect 207850 19410 208000 19480
rect 204000 19400 208000 19410
rect 204000 19380 204120 19400
rect 204380 19380 204620 19400
rect 204880 19380 205120 19400
rect 205380 19380 205620 19400
rect 205880 19380 206120 19400
rect 206380 19380 206620 19400
rect 206880 19380 207120 19400
rect 207380 19380 207620 19400
rect 207880 19380 208000 19400
rect 204000 19350 204100 19380
rect 204000 19150 204020 19350
rect 204090 19150 204100 19350
rect 204000 19120 204100 19150
rect 204400 19350 204600 19380
rect 204400 19150 204410 19350
rect 204480 19150 204520 19350
rect 204590 19150 204600 19350
rect 204400 19120 204600 19150
rect 204900 19350 205100 19380
rect 204900 19150 204910 19350
rect 204980 19150 205020 19350
rect 205090 19150 205100 19350
rect 204900 19120 205100 19150
rect 205400 19350 205600 19380
rect 205400 19150 205410 19350
rect 205480 19150 205520 19350
rect 205590 19150 205600 19350
rect 205400 19120 205600 19150
rect 205900 19350 206100 19380
rect 205900 19150 205910 19350
rect 205980 19150 206020 19350
rect 206090 19150 206100 19350
rect 205900 19120 206100 19150
rect 206400 19350 206600 19380
rect 206400 19150 206410 19350
rect 206480 19150 206520 19350
rect 206590 19150 206600 19350
rect 206400 19120 206600 19150
rect 206900 19350 207100 19380
rect 206900 19150 206910 19350
rect 206980 19150 207020 19350
rect 207090 19150 207100 19350
rect 206900 19120 207100 19150
rect 207400 19350 207600 19380
rect 207400 19150 207410 19350
rect 207480 19150 207520 19350
rect 207590 19150 207600 19350
rect 207400 19120 207600 19150
rect 207900 19350 208000 19380
rect 207900 19150 207910 19350
rect 207980 19150 208000 19350
rect 207900 19120 208000 19150
rect 204000 19100 204120 19120
rect 204380 19100 204620 19120
rect 204880 19100 205120 19120
rect 205380 19100 205620 19120
rect 205880 19100 206120 19120
rect 206380 19100 206620 19120
rect 206880 19100 207120 19120
rect 207380 19100 207620 19120
rect 207880 19100 208000 19120
rect 204000 19090 208000 19100
rect 204000 19020 204150 19090
rect 204350 19020 204650 19090
rect 204850 19020 205150 19090
rect 205350 19020 205650 19090
rect 205850 19020 206150 19090
rect 206350 19020 206650 19090
rect 206850 19020 207150 19090
rect 207350 19020 207650 19090
rect 207850 19020 208000 19090
rect 204000 18980 208000 19020
rect 204000 18910 204150 18980
rect 204350 18910 204650 18980
rect 204850 18910 205150 18980
rect 205350 18910 205650 18980
rect 205850 18910 206150 18980
rect 206350 18910 206650 18980
rect 206850 18910 207150 18980
rect 207350 18910 207650 18980
rect 207850 18910 208000 18980
rect 204000 18900 208000 18910
rect 204000 18880 204120 18900
rect 204380 18880 204620 18900
rect 204880 18880 205120 18900
rect 205380 18880 205620 18900
rect 205880 18880 206120 18900
rect 206380 18880 206620 18900
rect 206880 18880 207120 18900
rect 207380 18880 207620 18900
rect 207880 18880 208000 18900
rect 204000 18850 204100 18880
rect 204000 18650 204020 18850
rect 204090 18650 204100 18850
rect 204000 18620 204100 18650
rect 204400 18850 204600 18880
rect 204400 18650 204410 18850
rect 204480 18650 204520 18850
rect 204590 18650 204600 18850
rect 204400 18620 204600 18650
rect 204900 18850 205100 18880
rect 204900 18650 204910 18850
rect 204980 18650 205020 18850
rect 205090 18650 205100 18850
rect 204900 18620 205100 18650
rect 205400 18850 205600 18880
rect 205400 18650 205410 18850
rect 205480 18650 205520 18850
rect 205590 18650 205600 18850
rect 205400 18620 205600 18650
rect 205900 18850 206100 18880
rect 205900 18650 205910 18850
rect 205980 18650 206020 18850
rect 206090 18650 206100 18850
rect 205900 18620 206100 18650
rect 206400 18850 206600 18880
rect 206400 18650 206410 18850
rect 206480 18650 206520 18850
rect 206590 18650 206600 18850
rect 206400 18620 206600 18650
rect 206900 18850 207100 18880
rect 206900 18650 206910 18850
rect 206980 18650 207020 18850
rect 207090 18650 207100 18850
rect 206900 18620 207100 18650
rect 207400 18850 207600 18880
rect 207400 18650 207410 18850
rect 207480 18650 207520 18850
rect 207590 18650 207600 18850
rect 207400 18620 207600 18650
rect 207900 18850 208000 18880
rect 207900 18650 207910 18850
rect 207980 18650 208000 18850
rect 207900 18620 208000 18650
rect 204000 18600 204120 18620
rect 204380 18600 204620 18620
rect 204880 18600 205120 18620
rect 205380 18600 205620 18620
rect 205880 18600 206120 18620
rect 206380 18600 206620 18620
rect 206880 18600 207120 18620
rect 207380 18600 207620 18620
rect 207880 18600 208000 18620
rect 204000 18590 208000 18600
rect 204000 18520 204150 18590
rect 204350 18520 204650 18590
rect 204850 18520 205150 18590
rect 205350 18520 205650 18590
rect 205850 18520 206150 18590
rect 206350 18520 206650 18590
rect 206850 18520 207150 18590
rect 207350 18520 207650 18590
rect 207850 18520 208000 18590
rect 204000 18480 208000 18520
rect 204000 18410 204150 18480
rect 204350 18410 204650 18480
rect 204850 18410 205150 18480
rect 205350 18410 205650 18480
rect 205850 18410 206150 18480
rect 206350 18410 206650 18480
rect 206850 18410 207150 18480
rect 207350 18410 207650 18480
rect 207850 18410 208000 18480
rect 204000 18400 208000 18410
rect 204000 18380 204120 18400
rect 204380 18380 204620 18400
rect 204880 18380 205120 18400
rect 205380 18380 205620 18400
rect 205880 18380 206120 18400
rect 206380 18380 206620 18400
rect 206880 18380 207120 18400
rect 207380 18380 207620 18400
rect 207880 18380 208000 18400
rect 204000 18350 204100 18380
rect 204000 18150 204020 18350
rect 204090 18150 204100 18350
rect 204000 18120 204100 18150
rect 204400 18350 204600 18380
rect 204400 18150 204410 18350
rect 204480 18150 204520 18350
rect 204590 18150 204600 18350
rect 204400 18120 204600 18150
rect 204900 18350 205100 18380
rect 204900 18150 204910 18350
rect 204980 18150 205020 18350
rect 205090 18150 205100 18350
rect 204900 18120 205100 18150
rect 205400 18350 205600 18380
rect 205400 18150 205410 18350
rect 205480 18150 205520 18350
rect 205590 18150 205600 18350
rect 205400 18120 205600 18150
rect 205900 18350 206100 18380
rect 205900 18150 205910 18350
rect 205980 18150 206020 18350
rect 206090 18150 206100 18350
rect 205900 18120 206100 18150
rect 206400 18350 206600 18380
rect 206400 18150 206410 18350
rect 206480 18150 206520 18350
rect 206590 18150 206600 18350
rect 206400 18120 206600 18150
rect 206900 18350 207100 18380
rect 206900 18150 206910 18350
rect 206980 18150 207020 18350
rect 207090 18150 207100 18350
rect 206900 18120 207100 18150
rect 207400 18350 207600 18380
rect 207400 18150 207410 18350
rect 207480 18150 207520 18350
rect 207590 18150 207600 18350
rect 207400 18120 207600 18150
rect 207900 18350 208000 18380
rect 207900 18150 207910 18350
rect 207980 18150 208000 18350
rect 207900 18120 208000 18150
rect 204000 18100 204120 18120
rect 204380 18100 204620 18120
rect 204880 18100 205120 18120
rect 205380 18100 205620 18120
rect 205880 18100 206120 18120
rect 206380 18100 206620 18120
rect 206880 18100 207120 18120
rect 207380 18100 207620 18120
rect 207880 18100 208000 18120
rect 204000 18090 208000 18100
rect 204000 18020 204150 18090
rect 204350 18020 204650 18090
rect 204850 18020 205150 18090
rect 205350 18020 205650 18090
rect 205850 18020 206150 18090
rect 206350 18020 206650 18090
rect 206850 18020 207150 18090
rect 207350 18020 207650 18090
rect 207850 18020 208000 18090
rect 204000 17980 208000 18020
rect 204000 17910 204150 17980
rect 204350 17910 204650 17980
rect 204850 17910 205150 17980
rect 205350 17910 205650 17980
rect 205850 17910 206150 17980
rect 206350 17910 206650 17980
rect 206850 17910 207150 17980
rect 207350 17910 207650 17980
rect 207850 17910 208000 17980
rect 204000 17900 208000 17910
rect 204000 17880 204120 17900
rect 204380 17880 204620 17900
rect 204880 17880 205120 17900
rect 205380 17880 205620 17900
rect 205880 17880 206120 17900
rect 206380 17880 206620 17900
rect 206880 17880 207120 17900
rect 207380 17880 207620 17900
rect 207880 17880 208000 17900
rect 204000 17850 204100 17880
rect 204000 17650 204020 17850
rect 204090 17650 204100 17850
rect 204000 17620 204100 17650
rect 204400 17850 204600 17880
rect 204400 17650 204410 17850
rect 204480 17650 204520 17850
rect 204590 17650 204600 17850
rect 204400 17620 204600 17650
rect 204900 17850 205100 17880
rect 204900 17650 204910 17850
rect 204980 17650 205020 17850
rect 205090 17650 205100 17850
rect 204900 17620 205100 17650
rect 205400 17850 205600 17880
rect 205400 17650 205410 17850
rect 205480 17650 205520 17850
rect 205590 17650 205600 17850
rect 205400 17620 205600 17650
rect 205900 17850 206100 17880
rect 205900 17650 205910 17850
rect 205980 17650 206020 17850
rect 206090 17650 206100 17850
rect 205900 17620 206100 17650
rect 206400 17850 206600 17880
rect 206400 17650 206410 17850
rect 206480 17650 206520 17850
rect 206590 17650 206600 17850
rect 206400 17620 206600 17650
rect 206900 17850 207100 17880
rect 206900 17650 206910 17850
rect 206980 17650 207020 17850
rect 207090 17650 207100 17850
rect 206900 17620 207100 17650
rect 207400 17850 207600 17880
rect 207400 17650 207410 17850
rect 207480 17650 207520 17850
rect 207590 17650 207600 17850
rect 207400 17620 207600 17650
rect 207900 17850 208000 17880
rect 207900 17650 207910 17850
rect 207980 17650 208000 17850
rect 207900 17620 208000 17650
rect 204000 17600 204120 17620
rect 204380 17600 204620 17620
rect 204880 17600 205120 17620
rect 205380 17600 205620 17620
rect 205880 17600 206120 17620
rect 206380 17600 206620 17620
rect 206880 17600 207120 17620
rect 207380 17600 207620 17620
rect 207880 17600 208000 17620
rect 204000 17590 208000 17600
rect 204000 17520 204150 17590
rect 204350 17520 204650 17590
rect 204850 17520 205150 17590
rect 205350 17520 205650 17590
rect 205850 17520 206150 17590
rect 206350 17520 206650 17590
rect 206850 17520 207150 17590
rect 207350 17520 207650 17590
rect 207850 17520 208000 17590
rect 204000 17480 208000 17520
rect 204000 17410 204150 17480
rect 204350 17410 204650 17480
rect 204850 17410 205150 17480
rect 205350 17410 205650 17480
rect 205850 17410 206150 17480
rect 206350 17410 206650 17480
rect 206850 17410 207150 17480
rect 207350 17410 207650 17480
rect 207850 17410 208000 17480
rect 204000 17400 208000 17410
rect 204000 17380 204120 17400
rect 204380 17380 204620 17400
rect 204880 17380 205120 17400
rect 205380 17380 205620 17400
rect 205880 17380 206120 17400
rect 206380 17380 206620 17400
rect 206880 17380 207120 17400
rect 207380 17380 207620 17400
rect 207880 17380 208000 17400
rect 204000 17350 204100 17380
rect 204000 17150 204020 17350
rect 204090 17150 204100 17350
rect 204000 17120 204100 17150
rect 204400 17350 204600 17380
rect 204400 17150 204410 17350
rect 204480 17150 204520 17350
rect 204590 17150 204600 17350
rect 204400 17120 204600 17150
rect 204900 17350 205100 17380
rect 204900 17150 204910 17350
rect 204980 17150 205020 17350
rect 205090 17150 205100 17350
rect 204900 17120 205100 17150
rect 205400 17350 205600 17380
rect 205400 17150 205410 17350
rect 205480 17150 205520 17350
rect 205590 17150 205600 17350
rect 205400 17120 205600 17150
rect 205900 17350 206100 17380
rect 205900 17150 205910 17350
rect 205980 17150 206020 17350
rect 206090 17150 206100 17350
rect 205900 17120 206100 17150
rect 206400 17350 206600 17380
rect 206400 17150 206410 17350
rect 206480 17150 206520 17350
rect 206590 17150 206600 17350
rect 206400 17120 206600 17150
rect 206900 17350 207100 17380
rect 206900 17150 206910 17350
rect 206980 17150 207020 17350
rect 207090 17150 207100 17350
rect 206900 17120 207100 17150
rect 207400 17350 207600 17380
rect 207400 17150 207410 17350
rect 207480 17150 207520 17350
rect 207590 17150 207600 17350
rect 207400 17120 207600 17150
rect 207900 17350 208000 17380
rect 207900 17150 207910 17350
rect 207980 17150 208000 17350
rect 207900 17120 208000 17150
rect 204000 17100 204120 17120
rect 204380 17100 204620 17120
rect 204880 17100 205120 17120
rect 205380 17100 205620 17120
rect 205880 17100 206120 17120
rect 206380 17100 206620 17120
rect 206880 17100 207120 17120
rect 207380 17100 207620 17120
rect 207880 17100 208000 17120
rect 204000 17090 208000 17100
rect 204000 17020 204150 17090
rect 204350 17020 204650 17090
rect 204850 17020 205150 17090
rect 205350 17020 205650 17090
rect 205850 17020 206150 17090
rect 206350 17020 206650 17090
rect 206850 17020 207150 17090
rect 207350 17020 207650 17090
rect 207850 17020 208000 17090
rect 204000 16980 208000 17020
rect 204000 16910 204150 16980
rect 204350 16910 204650 16980
rect 204850 16910 205150 16980
rect 205350 16910 205650 16980
rect 205850 16910 206150 16980
rect 206350 16910 206650 16980
rect 206850 16910 207150 16980
rect 207350 16910 207650 16980
rect 207850 16910 208000 16980
rect 204000 16900 208000 16910
rect 204000 16880 204120 16900
rect 204380 16880 204620 16900
rect 204880 16880 205120 16900
rect 205380 16880 205620 16900
rect 205880 16880 206120 16900
rect 206380 16880 206620 16900
rect 206880 16880 207120 16900
rect 207380 16880 207620 16900
rect 207880 16880 208000 16900
rect 204000 16850 204100 16880
rect 204000 16650 204020 16850
rect 204090 16650 204100 16850
rect 204000 16620 204100 16650
rect 204400 16850 204600 16880
rect 204400 16650 204410 16850
rect 204480 16650 204520 16850
rect 204590 16650 204600 16850
rect 204400 16620 204600 16650
rect 204900 16850 205100 16880
rect 204900 16650 204910 16850
rect 204980 16650 205020 16850
rect 205090 16650 205100 16850
rect 204900 16620 205100 16650
rect 205400 16850 205600 16880
rect 205400 16650 205410 16850
rect 205480 16650 205520 16850
rect 205590 16650 205600 16850
rect 205400 16620 205600 16650
rect 205900 16850 206100 16880
rect 205900 16650 205910 16850
rect 205980 16650 206020 16850
rect 206090 16650 206100 16850
rect 205900 16620 206100 16650
rect 206400 16850 206600 16880
rect 206400 16650 206410 16850
rect 206480 16650 206520 16850
rect 206590 16650 206600 16850
rect 206400 16620 206600 16650
rect 206900 16850 207100 16880
rect 206900 16650 206910 16850
rect 206980 16650 207020 16850
rect 207090 16650 207100 16850
rect 206900 16620 207100 16650
rect 207400 16850 207600 16880
rect 207400 16650 207410 16850
rect 207480 16650 207520 16850
rect 207590 16650 207600 16850
rect 207400 16620 207600 16650
rect 207900 16850 208000 16880
rect 207900 16650 207910 16850
rect 207980 16650 208000 16850
rect 207900 16620 208000 16650
rect 204000 16600 204120 16620
rect 204380 16600 204620 16620
rect 204880 16600 205120 16620
rect 205380 16600 205620 16620
rect 205880 16600 206120 16620
rect 206380 16600 206620 16620
rect 206880 16600 207120 16620
rect 207380 16600 207620 16620
rect 207880 16600 208000 16620
rect 204000 16590 208000 16600
rect 204000 16520 204150 16590
rect 204350 16520 204650 16590
rect 204850 16520 205150 16590
rect 205350 16520 205650 16590
rect 205850 16520 206150 16590
rect 206350 16520 206650 16590
rect 206850 16520 207150 16590
rect 207350 16520 207650 16590
rect 207850 16520 208000 16590
rect 204000 16480 208000 16520
rect 204000 16410 204150 16480
rect 204350 16410 204650 16480
rect 204850 16410 205150 16480
rect 205350 16410 205650 16480
rect 205850 16410 206150 16480
rect 206350 16410 206650 16480
rect 206850 16410 207150 16480
rect 207350 16410 207650 16480
rect 207850 16410 208000 16480
rect 204000 16400 208000 16410
rect 204000 16380 204120 16400
rect 204380 16380 204620 16400
rect 204880 16380 205120 16400
rect 205380 16380 205620 16400
rect 205880 16380 206120 16400
rect 206380 16380 206620 16400
rect 206880 16380 207120 16400
rect 207380 16380 207620 16400
rect 207880 16380 208000 16400
rect 204000 16350 204100 16380
rect 204000 16150 204020 16350
rect 204090 16150 204100 16350
rect 204000 16120 204100 16150
rect 204400 16350 204600 16380
rect 204400 16150 204410 16350
rect 204480 16150 204520 16350
rect 204590 16150 204600 16350
rect 204400 16120 204600 16150
rect 204900 16350 205100 16380
rect 204900 16150 204910 16350
rect 204980 16150 205020 16350
rect 205090 16150 205100 16350
rect 204900 16120 205100 16150
rect 205400 16350 205600 16380
rect 205400 16150 205410 16350
rect 205480 16150 205520 16350
rect 205590 16150 205600 16350
rect 205400 16120 205600 16150
rect 205900 16350 206100 16380
rect 205900 16150 205910 16350
rect 205980 16150 206020 16350
rect 206090 16150 206100 16350
rect 205900 16120 206100 16150
rect 206400 16350 206600 16380
rect 206400 16150 206410 16350
rect 206480 16150 206520 16350
rect 206590 16150 206600 16350
rect 206400 16120 206600 16150
rect 206900 16350 207100 16380
rect 206900 16150 206910 16350
rect 206980 16150 207020 16350
rect 207090 16150 207100 16350
rect 206900 16120 207100 16150
rect 207400 16350 207600 16380
rect 207400 16150 207410 16350
rect 207480 16150 207520 16350
rect 207590 16150 207600 16350
rect 207400 16120 207600 16150
rect 207900 16350 208000 16380
rect 207900 16150 207910 16350
rect 207980 16150 208000 16350
rect 207900 16120 208000 16150
rect 204000 16100 204120 16120
rect 204380 16100 204620 16120
rect 204880 16100 205120 16120
rect 205380 16100 205620 16120
rect 205880 16100 206120 16120
rect 206380 16100 206620 16120
rect 206880 16100 207120 16120
rect 207380 16100 207620 16120
rect 207880 16100 208000 16120
rect 204000 16090 208000 16100
rect 204000 16020 204150 16090
rect 204350 16020 204650 16090
rect 204850 16020 205150 16090
rect 205350 16020 205650 16090
rect 205850 16020 206150 16090
rect 206350 16020 206650 16090
rect 206850 16020 207150 16090
rect 207350 16020 207650 16090
rect 207850 16020 208000 16090
rect 204000 15980 208000 16020
rect 204000 15910 204150 15980
rect 204350 15910 204650 15980
rect 204850 15910 205150 15980
rect 205350 15910 205650 15980
rect 205850 15910 206150 15980
rect 206350 15910 206650 15980
rect 206850 15910 207150 15980
rect 207350 15910 207650 15980
rect 207850 15910 208000 15980
rect 204000 15900 208000 15910
rect 204000 15880 204120 15900
rect 204380 15880 204620 15900
rect 204880 15880 205120 15900
rect 205380 15880 205620 15900
rect 205880 15880 206120 15900
rect 206380 15880 206620 15900
rect 206880 15880 207120 15900
rect 207380 15880 207620 15900
rect 207880 15880 208000 15900
rect 204000 15850 204100 15880
rect 204000 15650 204020 15850
rect 204090 15650 204100 15850
rect 204000 15620 204100 15650
rect 204400 15850 204600 15880
rect 204400 15650 204410 15850
rect 204480 15650 204520 15850
rect 204590 15650 204600 15850
rect 204400 15620 204600 15650
rect 204900 15850 205100 15880
rect 204900 15650 204910 15850
rect 204980 15650 205020 15850
rect 205090 15650 205100 15850
rect 204900 15620 205100 15650
rect 205400 15850 205600 15880
rect 205400 15650 205410 15850
rect 205480 15650 205520 15850
rect 205590 15650 205600 15850
rect 205400 15620 205600 15650
rect 205900 15850 206100 15880
rect 205900 15650 205910 15850
rect 205980 15650 206020 15850
rect 206090 15650 206100 15850
rect 205900 15620 206100 15650
rect 206400 15850 206600 15880
rect 206400 15650 206410 15850
rect 206480 15650 206520 15850
rect 206590 15650 206600 15850
rect 206400 15620 206600 15650
rect 206900 15850 207100 15880
rect 206900 15650 206910 15850
rect 206980 15650 207020 15850
rect 207090 15650 207100 15850
rect 206900 15620 207100 15650
rect 207400 15850 207600 15880
rect 207400 15650 207410 15850
rect 207480 15650 207520 15850
rect 207590 15650 207600 15850
rect 207400 15620 207600 15650
rect 207900 15850 208000 15880
rect 207900 15650 207910 15850
rect 207980 15650 208000 15850
rect 207900 15620 208000 15650
rect 204000 15600 204120 15620
rect 204380 15600 204620 15620
rect 204880 15600 205120 15620
rect 205380 15600 205620 15620
rect 205880 15600 206120 15620
rect 206380 15600 206620 15620
rect 206880 15600 207120 15620
rect 207380 15600 207620 15620
rect 207880 15600 208000 15620
rect 204000 15590 208000 15600
rect 204000 15520 204150 15590
rect 204350 15520 204650 15590
rect 204850 15520 205150 15590
rect 205350 15520 205650 15590
rect 205850 15520 206150 15590
rect 206350 15520 206650 15590
rect 206850 15520 207150 15590
rect 207350 15520 207650 15590
rect 207850 15520 208000 15590
rect 204000 15480 208000 15520
rect 204000 15410 204150 15480
rect 204350 15410 204650 15480
rect 204850 15410 205150 15480
rect 205350 15410 205650 15480
rect 205850 15410 206150 15480
rect 206350 15410 206650 15480
rect 206850 15410 207150 15480
rect 207350 15410 207650 15480
rect 207850 15410 208000 15480
rect 204000 15400 208000 15410
rect 204000 15380 204120 15400
rect 204380 15380 204620 15400
rect 204880 15380 205120 15400
rect 205380 15380 205620 15400
rect 205880 15380 206120 15400
rect 206380 15380 206620 15400
rect 206880 15380 207120 15400
rect 207380 15380 207620 15400
rect 207880 15380 208000 15400
rect 204000 15350 204100 15380
rect 204000 15150 204020 15350
rect 204090 15150 204100 15350
rect 204000 15120 204100 15150
rect 204400 15350 204600 15380
rect 204400 15150 204410 15350
rect 204480 15150 204520 15350
rect 204590 15150 204600 15350
rect 204400 15120 204600 15150
rect 204900 15350 205100 15380
rect 204900 15150 204910 15350
rect 204980 15150 205020 15350
rect 205090 15150 205100 15350
rect 204900 15120 205100 15150
rect 205400 15350 205600 15380
rect 205400 15150 205410 15350
rect 205480 15150 205520 15350
rect 205590 15150 205600 15350
rect 205400 15120 205600 15150
rect 205900 15350 206100 15380
rect 205900 15150 205910 15350
rect 205980 15150 206020 15350
rect 206090 15150 206100 15350
rect 205900 15120 206100 15150
rect 206400 15350 206600 15380
rect 206400 15150 206410 15350
rect 206480 15150 206520 15350
rect 206590 15150 206600 15350
rect 206400 15120 206600 15150
rect 206900 15350 207100 15380
rect 206900 15150 206910 15350
rect 206980 15150 207020 15350
rect 207090 15150 207100 15350
rect 206900 15120 207100 15150
rect 207400 15350 207600 15380
rect 207400 15150 207410 15350
rect 207480 15150 207520 15350
rect 207590 15150 207600 15350
rect 207400 15120 207600 15150
rect 207900 15350 208000 15380
rect 207900 15150 207910 15350
rect 207980 15150 208000 15350
rect 207900 15120 208000 15150
rect 204000 15100 204120 15120
rect 204380 15100 204620 15120
rect 204880 15100 205120 15120
rect 205380 15100 205620 15120
rect 205880 15100 206120 15120
rect 206380 15100 206620 15120
rect 206880 15100 207120 15120
rect 207380 15100 207620 15120
rect 207880 15100 208000 15120
rect 204000 15090 208000 15100
rect 204000 15020 204150 15090
rect 204350 15020 204650 15090
rect 204850 15020 205150 15090
rect 205350 15020 205650 15090
rect 205850 15020 206150 15090
rect 206350 15020 206650 15090
rect 206850 15020 207150 15090
rect 207350 15020 207650 15090
rect 207850 15020 208000 15090
rect 204000 14980 208000 15020
rect 204000 14910 204150 14980
rect 204350 14910 204650 14980
rect 204850 14910 205150 14980
rect 205350 14910 205650 14980
rect 205850 14910 206150 14980
rect 206350 14910 206650 14980
rect 206850 14910 207150 14980
rect 207350 14910 207650 14980
rect 207850 14910 208000 14980
rect 204000 14900 208000 14910
rect 204000 14880 204120 14900
rect 204380 14880 204620 14900
rect 204880 14880 205120 14900
rect 205380 14880 205620 14900
rect 205880 14880 206120 14900
rect 206380 14880 206620 14900
rect 206880 14880 207120 14900
rect 207380 14880 207620 14900
rect 207880 14880 208000 14900
rect 204000 14850 204100 14880
rect 204000 14650 204020 14850
rect 204090 14650 204100 14850
rect 204000 14620 204100 14650
rect 204400 14850 204600 14880
rect 204400 14650 204410 14850
rect 204480 14650 204520 14850
rect 204590 14650 204600 14850
rect 204400 14620 204600 14650
rect 204900 14850 205100 14880
rect 204900 14650 204910 14850
rect 204980 14650 205020 14850
rect 205090 14650 205100 14850
rect 204900 14620 205100 14650
rect 205400 14850 205600 14880
rect 205400 14650 205410 14850
rect 205480 14650 205520 14850
rect 205590 14650 205600 14850
rect 205400 14620 205600 14650
rect 205900 14850 206100 14880
rect 205900 14650 205910 14850
rect 205980 14650 206020 14850
rect 206090 14650 206100 14850
rect 205900 14620 206100 14650
rect 206400 14850 206600 14880
rect 206400 14650 206410 14850
rect 206480 14650 206520 14850
rect 206590 14650 206600 14850
rect 206400 14620 206600 14650
rect 206900 14850 207100 14880
rect 206900 14650 206910 14850
rect 206980 14650 207020 14850
rect 207090 14650 207100 14850
rect 206900 14620 207100 14650
rect 207400 14850 207600 14880
rect 207400 14650 207410 14850
rect 207480 14650 207520 14850
rect 207590 14650 207600 14850
rect 207400 14620 207600 14650
rect 207900 14850 208000 14880
rect 207900 14650 207910 14850
rect 207980 14650 208000 14850
rect 207900 14620 208000 14650
rect 204000 14600 204120 14620
rect 204380 14600 204620 14620
rect 204880 14600 205120 14620
rect 205380 14600 205620 14620
rect 205880 14600 206120 14620
rect 206380 14600 206620 14620
rect 206880 14600 207120 14620
rect 207380 14600 207620 14620
rect 207880 14600 208000 14620
rect 204000 14590 208000 14600
rect 204000 14520 204150 14590
rect 204350 14520 204650 14590
rect 204850 14520 205150 14590
rect 205350 14520 205650 14590
rect 205850 14520 206150 14590
rect 206350 14520 206650 14590
rect 206850 14520 207150 14590
rect 207350 14520 207650 14590
rect 207850 14520 208000 14590
rect 204000 14480 208000 14520
rect 204000 14410 204150 14480
rect 204350 14410 204650 14480
rect 204850 14410 205150 14480
rect 205350 14410 205650 14480
rect 205850 14410 206150 14480
rect 206350 14410 206650 14480
rect 206850 14410 207150 14480
rect 207350 14410 207650 14480
rect 207850 14410 208000 14480
rect 204000 14400 208000 14410
rect 204000 14380 204120 14400
rect 204380 14380 204620 14400
rect 204880 14380 205120 14400
rect 205380 14380 205620 14400
rect 205880 14380 206120 14400
rect 206380 14380 206620 14400
rect 206880 14380 207120 14400
rect 207380 14380 207620 14400
rect 207880 14380 208000 14400
rect 204000 14350 204100 14380
rect 204000 14150 204020 14350
rect 204090 14150 204100 14350
rect 204000 14120 204100 14150
rect 204400 14350 204600 14380
rect 204400 14150 204410 14350
rect 204480 14150 204520 14350
rect 204590 14150 204600 14350
rect 204400 14120 204600 14150
rect 204900 14350 205100 14380
rect 204900 14150 204910 14350
rect 204980 14150 205020 14350
rect 205090 14150 205100 14350
rect 204900 14120 205100 14150
rect 205400 14350 205600 14380
rect 205400 14150 205410 14350
rect 205480 14150 205520 14350
rect 205590 14150 205600 14350
rect 205400 14120 205600 14150
rect 205900 14350 206100 14380
rect 205900 14150 205910 14350
rect 205980 14150 206020 14350
rect 206090 14150 206100 14350
rect 205900 14120 206100 14150
rect 206400 14350 206600 14380
rect 206400 14150 206410 14350
rect 206480 14150 206520 14350
rect 206590 14150 206600 14350
rect 206400 14120 206600 14150
rect 206900 14350 207100 14380
rect 206900 14150 206910 14350
rect 206980 14150 207020 14350
rect 207090 14150 207100 14350
rect 206900 14120 207100 14150
rect 207400 14350 207600 14380
rect 207400 14150 207410 14350
rect 207480 14150 207520 14350
rect 207590 14150 207600 14350
rect 207400 14120 207600 14150
rect 207900 14350 208000 14380
rect 207900 14150 207910 14350
rect 207980 14150 208000 14350
rect 207900 14120 208000 14150
rect 204000 14100 204120 14120
rect 204380 14100 204620 14120
rect 204880 14100 205120 14120
rect 205380 14100 205620 14120
rect 205880 14100 206120 14120
rect 206380 14100 206620 14120
rect 206880 14100 207120 14120
rect 207380 14100 207620 14120
rect 207880 14100 208000 14120
rect 204000 14090 208000 14100
rect 204000 14020 204150 14090
rect 204350 14020 204650 14090
rect 204850 14020 205150 14090
rect 205350 14020 205650 14090
rect 205850 14020 206150 14090
rect 206350 14020 206650 14090
rect 206850 14020 207150 14090
rect 207350 14020 207650 14090
rect 207850 14020 208000 14090
rect 204000 13980 208000 14020
rect 204000 13910 204150 13980
rect 204350 13910 204650 13980
rect 204850 13910 205150 13980
rect 205350 13910 205650 13980
rect 205850 13910 206150 13980
rect 206350 13910 206650 13980
rect 206850 13910 207150 13980
rect 207350 13910 207650 13980
rect 207850 13910 208000 13980
rect 204000 13900 208000 13910
rect 204000 13880 204120 13900
rect 204380 13880 204620 13900
rect 204880 13880 205120 13900
rect 205380 13880 205620 13900
rect 205880 13880 206120 13900
rect 206380 13880 206620 13900
rect 206880 13880 207120 13900
rect 207380 13880 207620 13900
rect 207880 13880 208000 13900
rect 204000 13850 204100 13880
rect 204000 13650 204020 13850
rect 204090 13650 204100 13850
rect 204000 13620 204100 13650
rect 204400 13850 204600 13880
rect 204400 13650 204410 13850
rect 204480 13650 204520 13850
rect 204590 13650 204600 13850
rect 204400 13620 204600 13650
rect 204900 13850 205100 13880
rect 204900 13650 204910 13850
rect 204980 13650 205020 13850
rect 205090 13650 205100 13850
rect 204900 13620 205100 13650
rect 205400 13850 205600 13880
rect 205400 13650 205410 13850
rect 205480 13650 205520 13850
rect 205590 13650 205600 13850
rect 205400 13620 205600 13650
rect 205900 13850 206100 13880
rect 205900 13650 205910 13850
rect 205980 13650 206020 13850
rect 206090 13650 206100 13850
rect 205900 13620 206100 13650
rect 206400 13850 206600 13880
rect 206400 13650 206410 13850
rect 206480 13650 206520 13850
rect 206590 13650 206600 13850
rect 206400 13620 206600 13650
rect 206900 13850 207100 13880
rect 206900 13650 206910 13850
rect 206980 13650 207020 13850
rect 207090 13650 207100 13850
rect 206900 13620 207100 13650
rect 207400 13850 207600 13880
rect 207400 13650 207410 13850
rect 207480 13650 207520 13850
rect 207590 13650 207600 13850
rect 207400 13620 207600 13650
rect 207900 13850 208000 13880
rect 207900 13650 207910 13850
rect 207980 13650 208000 13850
rect 207900 13620 208000 13650
rect 204000 13600 204120 13620
rect 204380 13600 204620 13620
rect 204880 13600 205120 13620
rect 205380 13600 205620 13620
rect 205880 13600 206120 13620
rect 206380 13600 206620 13620
rect 206880 13600 207120 13620
rect 207380 13600 207620 13620
rect 207880 13600 208000 13620
rect 204000 13590 208000 13600
rect 204000 13520 204150 13590
rect 204350 13520 204650 13590
rect 204850 13520 205150 13590
rect 205350 13520 205650 13590
rect 205850 13520 206150 13590
rect 206350 13520 206650 13590
rect 206850 13520 207150 13590
rect 207350 13520 207650 13590
rect 207850 13520 208000 13590
rect 204000 13480 208000 13520
rect 204000 13410 204150 13480
rect 204350 13410 204650 13480
rect 204850 13410 205150 13480
rect 205350 13410 205650 13480
rect 205850 13410 206150 13480
rect 206350 13410 206650 13480
rect 206850 13410 207150 13480
rect 207350 13410 207650 13480
rect 207850 13410 208000 13480
rect 204000 13400 208000 13410
rect 204000 13380 204120 13400
rect 204380 13380 204620 13400
rect 204880 13380 205120 13400
rect 205380 13380 205620 13400
rect 205880 13380 206120 13400
rect 206380 13380 206620 13400
rect 206880 13380 207120 13400
rect 207380 13380 207620 13400
rect 207880 13380 208000 13400
rect 204000 13350 204100 13380
rect 204000 13150 204020 13350
rect 204090 13150 204100 13350
rect 204000 13120 204100 13150
rect 204400 13350 204600 13380
rect 204400 13150 204410 13350
rect 204480 13150 204520 13350
rect 204590 13150 204600 13350
rect 204400 13120 204600 13150
rect 204900 13350 205100 13380
rect 204900 13150 204910 13350
rect 204980 13150 205020 13350
rect 205090 13150 205100 13350
rect 204900 13120 205100 13150
rect 205400 13350 205600 13380
rect 205400 13150 205410 13350
rect 205480 13150 205520 13350
rect 205590 13150 205600 13350
rect 205400 13120 205600 13150
rect 205900 13350 206100 13380
rect 205900 13150 205910 13350
rect 205980 13150 206020 13350
rect 206090 13150 206100 13350
rect 205900 13120 206100 13150
rect 206400 13350 206600 13380
rect 206400 13150 206410 13350
rect 206480 13150 206520 13350
rect 206590 13150 206600 13350
rect 206400 13120 206600 13150
rect 206900 13350 207100 13380
rect 206900 13150 206910 13350
rect 206980 13150 207020 13350
rect 207090 13150 207100 13350
rect 206900 13120 207100 13150
rect 207400 13350 207600 13380
rect 207400 13150 207410 13350
rect 207480 13150 207520 13350
rect 207590 13150 207600 13350
rect 207400 13120 207600 13150
rect 207900 13350 208000 13380
rect 207900 13150 207910 13350
rect 207980 13150 208000 13350
rect 207900 13120 208000 13150
rect 204000 13100 204120 13120
rect 204380 13100 204620 13120
rect 204880 13100 205120 13120
rect 205380 13100 205620 13120
rect 205880 13100 206120 13120
rect 206380 13100 206620 13120
rect 206880 13100 207120 13120
rect 207380 13100 207620 13120
rect 207880 13100 208000 13120
rect 204000 13090 208000 13100
rect 204000 13020 204150 13090
rect 204350 13020 204650 13090
rect 204850 13020 205150 13090
rect 205350 13020 205650 13090
rect 205850 13020 206150 13090
rect 206350 13020 206650 13090
rect 206850 13020 207150 13090
rect 207350 13020 207650 13090
rect 207850 13020 208000 13090
rect 204000 12980 208000 13020
rect 204000 12910 204150 12980
rect 204350 12910 204650 12980
rect 204850 12910 205150 12980
rect 205350 12910 205650 12980
rect 205850 12910 206150 12980
rect 206350 12910 206650 12980
rect 206850 12910 207150 12980
rect 207350 12910 207650 12980
rect 207850 12910 208000 12980
rect 204000 12900 208000 12910
rect 204000 12880 204120 12900
rect 204380 12880 204620 12900
rect 204880 12880 205120 12900
rect 205380 12880 205620 12900
rect 205880 12880 206120 12900
rect 206380 12880 206620 12900
rect 206880 12880 207120 12900
rect 207380 12880 207620 12900
rect 207880 12880 208000 12900
rect 204000 12850 204100 12880
rect 204000 12650 204020 12850
rect 204090 12650 204100 12850
rect 204000 12620 204100 12650
rect 204400 12850 204600 12880
rect 204400 12650 204410 12850
rect 204480 12650 204520 12850
rect 204590 12650 204600 12850
rect 204400 12620 204600 12650
rect 204900 12850 205100 12880
rect 204900 12650 204910 12850
rect 204980 12650 205020 12850
rect 205090 12650 205100 12850
rect 204900 12620 205100 12650
rect 205400 12850 205600 12880
rect 205400 12650 205410 12850
rect 205480 12650 205520 12850
rect 205590 12650 205600 12850
rect 205400 12620 205600 12650
rect 205900 12850 206100 12880
rect 205900 12650 205910 12850
rect 205980 12650 206020 12850
rect 206090 12650 206100 12850
rect 205900 12620 206100 12650
rect 206400 12850 206600 12880
rect 206400 12650 206410 12850
rect 206480 12650 206520 12850
rect 206590 12650 206600 12850
rect 206400 12620 206600 12650
rect 206900 12850 207100 12880
rect 206900 12650 206910 12850
rect 206980 12650 207020 12850
rect 207090 12650 207100 12850
rect 206900 12620 207100 12650
rect 207400 12850 207600 12880
rect 207400 12650 207410 12850
rect 207480 12650 207520 12850
rect 207590 12650 207600 12850
rect 207400 12620 207600 12650
rect 207900 12850 208000 12880
rect 207900 12650 207910 12850
rect 207980 12650 208000 12850
rect 207900 12620 208000 12650
rect 204000 12600 204120 12620
rect 204380 12600 204620 12620
rect 204880 12600 205120 12620
rect 205380 12600 205620 12620
rect 205880 12600 206120 12620
rect 206380 12600 206620 12620
rect 206880 12600 207120 12620
rect 207380 12600 207620 12620
rect 207880 12600 208000 12620
rect 204000 12590 208000 12600
rect 204000 12520 204150 12590
rect 204350 12520 204650 12590
rect 204850 12520 205150 12590
rect 205350 12520 205650 12590
rect 205850 12520 206150 12590
rect 206350 12520 206650 12590
rect 206850 12520 207150 12590
rect 207350 12520 207650 12590
rect 207850 12520 208000 12590
rect 204000 12480 208000 12520
rect 204000 12410 204150 12480
rect 204350 12410 204650 12480
rect 204850 12410 205150 12480
rect 205350 12410 205650 12480
rect 205850 12410 206150 12480
rect 206350 12410 206650 12480
rect 206850 12410 207150 12480
rect 207350 12410 207650 12480
rect 207850 12410 208000 12480
rect 204000 12400 208000 12410
rect 204000 12380 204120 12400
rect 204380 12380 204620 12400
rect 204880 12380 205120 12400
rect 205380 12380 205620 12400
rect 205880 12380 206120 12400
rect 206380 12380 206620 12400
rect 206880 12380 207120 12400
rect 207380 12380 207620 12400
rect 207880 12380 208000 12400
rect 204000 12350 204100 12380
rect 204000 12150 204020 12350
rect 204090 12150 204100 12350
rect 204000 12120 204100 12150
rect 204400 12350 204600 12380
rect 204400 12150 204410 12350
rect 204480 12150 204520 12350
rect 204590 12150 204600 12350
rect 204400 12120 204600 12150
rect 204900 12350 205100 12380
rect 204900 12150 204910 12350
rect 204980 12150 205020 12350
rect 205090 12150 205100 12350
rect 204900 12120 205100 12150
rect 205400 12350 205600 12380
rect 205400 12150 205410 12350
rect 205480 12150 205520 12350
rect 205590 12150 205600 12350
rect 205400 12120 205600 12150
rect 205900 12350 206100 12380
rect 205900 12150 205910 12350
rect 205980 12150 206020 12350
rect 206090 12150 206100 12350
rect 205900 12120 206100 12150
rect 206400 12350 206600 12380
rect 206400 12150 206410 12350
rect 206480 12150 206520 12350
rect 206590 12150 206600 12350
rect 206400 12120 206600 12150
rect 206900 12350 207100 12380
rect 206900 12150 206910 12350
rect 206980 12150 207020 12350
rect 207090 12150 207100 12350
rect 206900 12120 207100 12150
rect 207400 12350 207600 12380
rect 207400 12150 207410 12350
rect 207480 12150 207520 12350
rect 207590 12150 207600 12350
rect 207400 12120 207600 12150
rect 207900 12350 208000 12380
rect 207900 12150 207910 12350
rect 207980 12150 208000 12350
rect 207900 12120 208000 12150
rect 204000 12100 204120 12120
rect 204380 12100 204620 12120
rect 204880 12100 205120 12120
rect 205380 12100 205620 12120
rect 205880 12100 206120 12120
rect 206380 12100 206620 12120
rect 206880 12100 207120 12120
rect 207380 12100 207620 12120
rect 207880 12100 208000 12120
rect 204000 12090 208000 12100
rect 204000 12020 204150 12090
rect 204350 12020 204650 12090
rect 204850 12020 205150 12090
rect 205350 12020 205650 12090
rect 205850 12020 206150 12090
rect 206350 12020 206650 12090
rect 206850 12020 207150 12090
rect 207350 12020 207650 12090
rect 207850 12020 208000 12090
rect 204000 11980 208000 12020
rect 204000 11910 204150 11980
rect 204350 11910 204650 11980
rect 204850 11910 205150 11980
rect 205350 11910 205650 11980
rect 205850 11910 206150 11980
rect 206350 11910 206650 11980
rect 206850 11910 207150 11980
rect 207350 11910 207650 11980
rect 207850 11910 208000 11980
rect 204000 11900 208000 11910
rect 204000 11880 204120 11900
rect 204380 11880 204620 11900
rect 204880 11880 205120 11900
rect 205380 11880 205620 11900
rect 205880 11880 206120 11900
rect 206380 11880 206620 11900
rect 206880 11880 207120 11900
rect 207380 11880 207620 11900
rect 207880 11880 208000 11900
rect 204000 11850 204100 11880
rect 204000 11650 204020 11850
rect 204090 11650 204100 11850
rect 204000 11620 204100 11650
rect 204400 11850 204600 11880
rect 204400 11650 204410 11850
rect 204480 11650 204520 11850
rect 204590 11650 204600 11850
rect 204400 11620 204600 11650
rect 204900 11850 205100 11880
rect 204900 11650 204910 11850
rect 204980 11650 205020 11850
rect 205090 11650 205100 11850
rect 204900 11620 205100 11650
rect 205400 11850 205600 11880
rect 205400 11650 205410 11850
rect 205480 11650 205520 11850
rect 205590 11650 205600 11850
rect 205400 11620 205600 11650
rect 205900 11850 206100 11880
rect 205900 11650 205910 11850
rect 205980 11650 206020 11850
rect 206090 11650 206100 11850
rect 205900 11620 206100 11650
rect 206400 11850 206600 11880
rect 206400 11650 206410 11850
rect 206480 11650 206520 11850
rect 206590 11650 206600 11850
rect 206400 11620 206600 11650
rect 206900 11850 207100 11880
rect 206900 11650 206910 11850
rect 206980 11650 207020 11850
rect 207090 11650 207100 11850
rect 206900 11620 207100 11650
rect 207400 11850 207600 11880
rect 207400 11650 207410 11850
rect 207480 11650 207520 11850
rect 207590 11650 207600 11850
rect 207400 11620 207600 11650
rect 207900 11850 208000 11880
rect 207900 11650 207910 11850
rect 207980 11650 208000 11850
rect 207900 11620 208000 11650
rect 204000 11600 204120 11620
rect 204380 11600 204620 11620
rect 204880 11600 205120 11620
rect 205380 11600 205620 11620
rect 205880 11600 206120 11620
rect 206380 11600 206620 11620
rect 206880 11600 207120 11620
rect 207380 11600 207620 11620
rect 207880 11600 208000 11620
rect 204000 11590 208000 11600
rect 204000 11520 204150 11590
rect 204350 11520 204650 11590
rect 204850 11520 205150 11590
rect 205350 11520 205650 11590
rect 205850 11520 206150 11590
rect 206350 11520 206650 11590
rect 206850 11520 207150 11590
rect 207350 11520 207650 11590
rect 207850 11520 208000 11590
rect 204000 11480 208000 11520
rect 204000 11410 204150 11480
rect 204350 11410 204650 11480
rect 204850 11410 205150 11480
rect 205350 11410 205650 11480
rect 205850 11410 206150 11480
rect 206350 11410 206650 11480
rect 206850 11410 207150 11480
rect 207350 11410 207650 11480
rect 207850 11410 208000 11480
rect 204000 11400 208000 11410
rect 204000 11380 204120 11400
rect 204380 11380 204620 11400
rect 204880 11380 205120 11400
rect 205380 11380 205620 11400
rect 205880 11380 206120 11400
rect 206380 11380 206620 11400
rect 206880 11380 207120 11400
rect 207380 11380 207620 11400
rect 207880 11380 208000 11400
rect 204000 11350 204100 11380
rect 204000 11150 204020 11350
rect 204090 11150 204100 11350
rect 204000 11120 204100 11150
rect 204400 11350 204600 11380
rect 204400 11150 204410 11350
rect 204480 11150 204520 11350
rect 204590 11150 204600 11350
rect 204400 11120 204600 11150
rect 204900 11350 205100 11380
rect 204900 11150 204910 11350
rect 204980 11150 205020 11350
rect 205090 11150 205100 11350
rect 204900 11120 205100 11150
rect 205400 11350 205600 11380
rect 205400 11150 205410 11350
rect 205480 11150 205520 11350
rect 205590 11150 205600 11350
rect 205400 11120 205600 11150
rect 205900 11350 206100 11380
rect 205900 11150 205910 11350
rect 205980 11150 206020 11350
rect 206090 11150 206100 11350
rect 205900 11120 206100 11150
rect 206400 11350 206600 11380
rect 206400 11150 206410 11350
rect 206480 11150 206520 11350
rect 206590 11150 206600 11350
rect 206400 11120 206600 11150
rect 206900 11350 207100 11380
rect 206900 11150 206910 11350
rect 206980 11150 207020 11350
rect 207090 11150 207100 11350
rect 206900 11120 207100 11150
rect 207400 11350 207600 11380
rect 207400 11150 207410 11350
rect 207480 11150 207520 11350
rect 207590 11150 207600 11350
rect 207400 11120 207600 11150
rect 207900 11350 208000 11380
rect 207900 11150 207910 11350
rect 207980 11150 208000 11350
rect 207900 11120 208000 11150
rect 204000 11100 204120 11120
rect 204380 11100 204620 11120
rect 204880 11100 205120 11120
rect 205380 11100 205620 11120
rect 205880 11100 206120 11120
rect 206380 11100 206620 11120
rect 206880 11100 207120 11120
rect 207380 11100 207620 11120
rect 207880 11100 208000 11120
rect 204000 11090 208000 11100
rect 204000 11020 204150 11090
rect 204350 11020 204650 11090
rect 204850 11020 205150 11090
rect 205350 11020 205650 11090
rect 205850 11020 206150 11090
rect 206350 11020 206650 11090
rect 206850 11020 207150 11090
rect 207350 11020 207650 11090
rect 207850 11020 208000 11090
rect 204000 10980 208000 11020
rect 204000 10910 204150 10980
rect 204350 10910 204650 10980
rect 204850 10910 205150 10980
rect 205350 10910 205650 10980
rect 205850 10910 206150 10980
rect 206350 10910 206650 10980
rect 206850 10910 207150 10980
rect 207350 10910 207650 10980
rect 207850 10910 208000 10980
rect 204000 10900 208000 10910
rect 204000 10880 204120 10900
rect 204380 10880 204620 10900
rect 204880 10880 205120 10900
rect 205380 10880 205620 10900
rect 205880 10880 206120 10900
rect 206380 10880 206620 10900
rect 206880 10880 207120 10900
rect 207380 10880 207620 10900
rect 207880 10880 208000 10900
rect 204000 10850 204100 10880
rect 204000 10650 204020 10850
rect 204090 10650 204100 10850
rect 204000 10620 204100 10650
rect 204400 10850 204600 10880
rect 204400 10650 204410 10850
rect 204480 10650 204520 10850
rect 204590 10650 204600 10850
rect 204400 10620 204600 10650
rect 204900 10850 205100 10880
rect 204900 10650 204910 10850
rect 204980 10650 205020 10850
rect 205090 10650 205100 10850
rect 204900 10620 205100 10650
rect 205400 10850 205600 10880
rect 205400 10650 205410 10850
rect 205480 10650 205520 10850
rect 205590 10650 205600 10850
rect 205400 10620 205600 10650
rect 205900 10850 206100 10880
rect 205900 10650 205910 10850
rect 205980 10650 206020 10850
rect 206090 10650 206100 10850
rect 205900 10620 206100 10650
rect 206400 10850 206600 10880
rect 206400 10650 206410 10850
rect 206480 10650 206520 10850
rect 206590 10650 206600 10850
rect 206400 10620 206600 10650
rect 206900 10850 207100 10880
rect 206900 10650 206910 10850
rect 206980 10650 207020 10850
rect 207090 10650 207100 10850
rect 206900 10620 207100 10650
rect 207400 10850 207600 10880
rect 207400 10650 207410 10850
rect 207480 10650 207520 10850
rect 207590 10650 207600 10850
rect 207400 10620 207600 10650
rect 207900 10850 208000 10880
rect 207900 10650 207910 10850
rect 207980 10650 208000 10850
rect 207900 10620 208000 10650
rect 204000 10600 204120 10620
rect 204380 10600 204620 10620
rect 204880 10600 205120 10620
rect 205380 10600 205620 10620
rect 205880 10600 206120 10620
rect 206380 10600 206620 10620
rect 206880 10600 207120 10620
rect 207380 10600 207620 10620
rect 207880 10600 208000 10620
rect 204000 10590 208000 10600
rect 204000 10520 204150 10590
rect 204350 10520 204650 10590
rect 204850 10520 205150 10590
rect 205350 10520 205650 10590
rect 205850 10520 206150 10590
rect 206350 10520 206650 10590
rect 206850 10520 207150 10590
rect 207350 10520 207650 10590
rect 207850 10520 208000 10590
rect 204000 10480 208000 10520
rect 204000 10410 204150 10480
rect 204350 10410 204650 10480
rect 204850 10410 205150 10480
rect 205350 10410 205650 10480
rect 205850 10410 206150 10480
rect 206350 10410 206650 10480
rect 206850 10410 207150 10480
rect 207350 10410 207650 10480
rect 207850 10410 208000 10480
rect 204000 10400 208000 10410
rect 204000 10380 204120 10400
rect 204380 10380 204620 10400
rect 204880 10380 205120 10400
rect 205380 10380 205620 10400
rect 205880 10380 206120 10400
rect 206380 10380 206620 10400
rect 206880 10380 207120 10400
rect 207380 10380 207620 10400
rect 207880 10380 208000 10400
rect 204000 10350 204100 10380
rect 204000 10150 204020 10350
rect 204090 10150 204100 10350
rect 204000 10120 204100 10150
rect 204400 10350 204600 10380
rect 204400 10150 204410 10350
rect 204480 10150 204520 10350
rect 204590 10150 204600 10350
rect 204400 10120 204600 10150
rect 204900 10350 205100 10380
rect 204900 10150 204910 10350
rect 204980 10150 205020 10350
rect 205090 10150 205100 10350
rect 204900 10120 205100 10150
rect 205400 10350 205600 10380
rect 205400 10150 205410 10350
rect 205480 10150 205520 10350
rect 205590 10150 205600 10350
rect 205400 10120 205600 10150
rect 205900 10350 206100 10380
rect 205900 10150 205910 10350
rect 205980 10150 206020 10350
rect 206090 10150 206100 10350
rect 205900 10120 206100 10150
rect 206400 10350 206600 10380
rect 206400 10150 206410 10350
rect 206480 10150 206520 10350
rect 206590 10150 206600 10350
rect 206400 10120 206600 10150
rect 206900 10350 207100 10380
rect 206900 10150 206910 10350
rect 206980 10150 207020 10350
rect 207090 10150 207100 10350
rect 206900 10120 207100 10150
rect 207400 10350 207600 10380
rect 207400 10150 207410 10350
rect 207480 10150 207520 10350
rect 207590 10150 207600 10350
rect 207400 10120 207600 10150
rect 207900 10350 208000 10380
rect 207900 10150 207910 10350
rect 207980 10150 208000 10350
rect 207900 10120 208000 10150
rect 204000 10100 204120 10120
rect 204380 10100 204620 10120
rect 204880 10100 205120 10120
rect 205380 10100 205620 10120
rect 205880 10100 206120 10120
rect 206380 10100 206620 10120
rect 206880 10100 207120 10120
rect 207380 10100 207620 10120
rect 207880 10100 208000 10120
rect 204000 10090 208000 10100
rect 204000 10020 204150 10090
rect 204350 10020 204650 10090
rect 204850 10020 205150 10090
rect 205350 10020 205650 10090
rect 205850 10020 206150 10090
rect 206350 10020 206650 10090
rect 206850 10020 207150 10090
rect 207350 10020 207650 10090
rect 207850 10020 208000 10090
rect 204000 9980 208000 10020
rect 204000 9910 204150 9980
rect 204350 9910 204650 9980
rect 204850 9910 205150 9980
rect 205350 9910 205650 9980
rect 205850 9910 206150 9980
rect 206350 9910 206650 9980
rect 206850 9910 207150 9980
rect 207350 9910 207650 9980
rect 207850 9910 208000 9980
rect 204000 9900 208000 9910
rect 204000 9880 204120 9900
rect 204380 9880 204620 9900
rect 204880 9880 205120 9900
rect 205380 9880 205620 9900
rect 205880 9880 206120 9900
rect 206380 9880 206620 9900
rect 206880 9880 207120 9900
rect 207380 9880 207620 9900
rect 207880 9880 208000 9900
rect 204000 9850 204100 9880
rect 204000 9650 204020 9850
rect 204090 9650 204100 9850
rect 204000 9620 204100 9650
rect 204400 9850 204600 9880
rect 204400 9650 204410 9850
rect 204480 9650 204520 9850
rect 204590 9650 204600 9850
rect 204400 9620 204600 9650
rect 204900 9850 205100 9880
rect 204900 9650 204910 9850
rect 204980 9650 205020 9850
rect 205090 9650 205100 9850
rect 204900 9620 205100 9650
rect 205400 9850 205600 9880
rect 205400 9650 205410 9850
rect 205480 9650 205520 9850
rect 205590 9650 205600 9850
rect 205400 9620 205600 9650
rect 205900 9850 206100 9880
rect 205900 9650 205910 9850
rect 205980 9650 206020 9850
rect 206090 9650 206100 9850
rect 205900 9620 206100 9650
rect 206400 9850 206600 9880
rect 206400 9650 206410 9850
rect 206480 9650 206520 9850
rect 206590 9650 206600 9850
rect 206400 9620 206600 9650
rect 206900 9850 207100 9880
rect 206900 9650 206910 9850
rect 206980 9650 207020 9850
rect 207090 9650 207100 9850
rect 206900 9620 207100 9650
rect 207400 9850 207600 9880
rect 207400 9650 207410 9850
rect 207480 9650 207520 9850
rect 207590 9650 207600 9850
rect 207400 9620 207600 9650
rect 207900 9850 208000 9880
rect 207900 9650 207910 9850
rect 207980 9650 208000 9850
rect 207900 9620 208000 9650
rect 204000 9600 204120 9620
rect 204380 9600 204620 9620
rect 204880 9600 205120 9620
rect 205380 9600 205620 9620
rect 205880 9600 206120 9620
rect 206380 9600 206620 9620
rect 206880 9600 207120 9620
rect 207380 9600 207620 9620
rect 207880 9600 208000 9620
rect 204000 9590 208000 9600
rect 204000 9520 204150 9590
rect 204350 9520 204650 9590
rect 204850 9520 205150 9590
rect 205350 9520 205650 9590
rect 205850 9520 206150 9590
rect 206350 9520 206650 9590
rect 206850 9520 207150 9590
rect 207350 9520 207650 9590
rect 207850 9520 208000 9590
rect 204000 9480 208000 9520
rect 204000 9410 204150 9480
rect 204350 9410 204650 9480
rect 204850 9410 205150 9480
rect 205350 9410 205650 9480
rect 205850 9410 206150 9480
rect 206350 9410 206650 9480
rect 206850 9410 207150 9480
rect 207350 9410 207650 9480
rect 207850 9410 208000 9480
rect 204000 9400 208000 9410
rect 204000 9380 204120 9400
rect 204380 9380 204620 9400
rect 204880 9380 205120 9400
rect 205380 9380 205620 9400
rect 205880 9380 206120 9400
rect 206380 9380 206620 9400
rect 206880 9380 207120 9400
rect 207380 9380 207620 9400
rect 207880 9380 208000 9400
rect 204000 9350 204100 9380
rect 204000 9150 204020 9350
rect 204090 9150 204100 9350
rect 204000 9120 204100 9150
rect 204400 9350 204600 9380
rect 204400 9150 204410 9350
rect 204480 9150 204520 9350
rect 204590 9150 204600 9350
rect 204400 9120 204600 9150
rect 204900 9350 205100 9380
rect 204900 9150 204910 9350
rect 204980 9150 205020 9350
rect 205090 9150 205100 9350
rect 204900 9120 205100 9150
rect 205400 9350 205600 9380
rect 205400 9150 205410 9350
rect 205480 9150 205520 9350
rect 205590 9150 205600 9350
rect 205400 9120 205600 9150
rect 205900 9350 206100 9380
rect 205900 9150 205910 9350
rect 205980 9150 206020 9350
rect 206090 9150 206100 9350
rect 205900 9120 206100 9150
rect 206400 9350 206600 9380
rect 206400 9150 206410 9350
rect 206480 9150 206520 9350
rect 206590 9150 206600 9350
rect 206400 9120 206600 9150
rect 206900 9350 207100 9380
rect 206900 9150 206910 9350
rect 206980 9150 207020 9350
rect 207090 9150 207100 9350
rect 206900 9120 207100 9150
rect 207400 9350 207600 9380
rect 207400 9150 207410 9350
rect 207480 9150 207520 9350
rect 207590 9150 207600 9350
rect 207400 9120 207600 9150
rect 207900 9350 208000 9380
rect 207900 9150 207910 9350
rect 207980 9150 208000 9350
rect 207900 9120 208000 9150
rect 204000 9100 204120 9120
rect 204380 9100 204620 9120
rect 204880 9100 205120 9120
rect 205380 9100 205620 9120
rect 205880 9100 206120 9120
rect 206380 9100 206620 9120
rect 206880 9100 207120 9120
rect 207380 9100 207620 9120
rect 207880 9100 208000 9120
rect 204000 9090 208000 9100
rect 204000 9020 204150 9090
rect 204350 9020 204650 9090
rect 204850 9020 205150 9090
rect 205350 9020 205650 9090
rect 205850 9020 206150 9090
rect 206350 9020 206650 9090
rect 206850 9020 207150 9090
rect 207350 9020 207650 9090
rect 207850 9020 208000 9090
rect 204000 8980 208000 9020
rect 204000 8910 204150 8980
rect 204350 8910 204650 8980
rect 204850 8910 205150 8980
rect 205350 8910 205650 8980
rect 205850 8910 206150 8980
rect 206350 8910 206650 8980
rect 206850 8910 207150 8980
rect 207350 8910 207650 8980
rect 207850 8910 208000 8980
rect 204000 8900 208000 8910
rect 204000 8880 204120 8900
rect 204380 8880 204620 8900
rect 204880 8880 205120 8900
rect 205380 8880 205620 8900
rect 205880 8880 206120 8900
rect 206380 8880 206620 8900
rect 206880 8880 207120 8900
rect 207380 8880 207620 8900
rect 207880 8880 208000 8900
rect 204000 8850 204100 8880
rect 204000 8650 204020 8850
rect 204090 8650 204100 8850
rect 204000 8620 204100 8650
rect 204400 8850 204600 8880
rect 204400 8650 204410 8850
rect 204480 8650 204520 8850
rect 204590 8650 204600 8850
rect 204400 8620 204600 8650
rect 204900 8850 205100 8880
rect 204900 8650 204910 8850
rect 204980 8650 205020 8850
rect 205090 8650 205100 8850
rect 204900 8620 205100 8650
rect 205400 8850 205600 8880
rect 205400 8650 205410 8850
rect 205480 8650 205520 8850
rect 205590 8650 205600 8850
rect 205400 8620 205600 8650
rect 205900 8850 206100 8880
rect 205900 8650 205910 8850
rect 205980 8650 206020 8850
rect 206090 8650 206100 8850
rect 205900 8620 206100 8650
rect 206400 8850 206600 8880
rect 206400 8650 206410 8850
rect 206480 8650 206520 8850
rect 206590 8650 206600 8850
rect 206400 8620 206600 8650
rect 206900 8850 207100 8880
rect 206900 8650 206910 8850
rect 206980 8650 207020 8850
rect 207090 8650 207100 8850
rect 206900 8620 207100 8650
rect 207400 8850 207600 8880
rect 207400 8650 207410 8850
rect 207480 8650 207520 8850
rect 207590 8650 207600 8850
rect 207400 8620 207600 8650
rect 207900 8850 208000 8880
rect 207900 8650 207910 8850
rect 207980 8650 208000 8850
rect 207900 8620 208000 8650
rect 204000 8600 204120 8620
rect 204380 8600 204620 8620
rect 204880 8600 205120 8620
rect 205380 8600 205620 8620
rect 205880 8600 206120 8620
rect 206380 8600 206620 8620
rect 206880 8600 207120 8620
rect 207380 8600 207620 8620
rect 207880 8600 208000 8620
rect 204000 8590 208000 8600
rect 204000 8520 204150 8590
rect 204350 8520 204650 8590
rect 204850 8520 205150 8590
rect 205350 8520 205650 8590
rect 205850 8520 206150 8590
rect 206350 8520 206650 8590
rect 206850 8520 207150 8590
rect 207350 8520 207650 8590
rect 207850 8520 208000 8590
rect 204000 8480 208000 8520
rect 204000 8410 204150 8480
rect 204350 8410 204650 8480
rect 204850 8410 205150 8480
rect 205350 8410 205650 8480
rect 205850 8410 206150 8480
rect 206350 8410 206650 8480
rect 206850 8410 207150 8480
rect 207350 8410 207650 8480
rect 207850 8410 208000 8480
rect 204000 8400 208000 8410
rect 204000 8380 204120 8400
rect 204380 8380 204620 8400
rect 204880 8380 205120 8400
rect 205380 8380 205620 8400
rect 205880 8380 206120 8400
rect 206380 8380 206620 8400
rect 206880 8380 207120 8400
rect 207380 8380 207620 8400
rect 207880 8380 208000 8400
rect 204000 8350 204100 8380
rect 204000 8150 204020 8350
rect 204090 8150 204100 8350
rect 204000 8120 204100 8150
rect 204400 8350 204600 8380
rect 204400 8150 204410 8350
rect 204480 8150 204520 8350
rect 204590 8150 204600 8350
rect 204400 8120 204600 8150
rect 204900 8350 205100 8380
rect 204900 8150 204910 8350
rect 204980 8150 205020 8350
rect 205090 8150 205100 8350
rect 204900 8120 205100 8150
rect 205400 8350 205600 8380
rect 205400 8150 205410 8350
rect 205480 8150 205520 8350
rect 205590 8150 205600 8350
rect 205400 8120 205600 8150
rect 205900 8350 206100 8380
rect 205900 8150 205910 8350
rect 205980 8150 206020 8350
rect 206090 8150 206100 8350
rect 205900 8120 206100 8150
rect 206400 8350 206600 8380
rect 206400 8150 206410 8350
rect 206480 8150 206520 8350
rect 206590 8150 206600 8350
rect 206400 8120 206600 8150
rect 206900 8350 207100 8380
rect 206900 8150 206910 8350
rect 206980 8150 207020 8350
rect 207090 8150 207100 8350
rect 206900 8120 207100 8150
rect 207400 8350 207600 8380
rect 207400 8150 207410 8350
rect 207480 8150 207520 8350
rect 207590 8150 207600 8350
rect 207400 8120 207600 8150
rect 207900 8350 208000 8380
rect 207900 8150 207910 8350
rect 207980 8150 208000 8350
rect 207900 8120 208000 8150
rect 204000 8100 204120 8120
rect 204380 8100 204620 8120
rect 204880 8100 205120 8120
rect 205380 8100 205620 8120
rect 205880 8100 206120 8120
rect 206380 8100 206620 8120
rect 206880 8100 207120 8120
rect 207380 8100 207620 8120
rect 207880 8100 208000 8120
rect 204000 8090 208000 8100
rect 204000 8020 204150 8090
rect 204350 8020 204650 8090
rect 204850 8020 205150 8090
rect 205350 8020 205650 8090
rect 205850 8020 206150 8090
rect 206350 8020 206650 8090
rect 206850 8020 207150 8090
rect 207350 8020 207650 8090
rect 207850 8020 208000 8090
rect 204000 7980 208000 8020
rect 204000 7910 204150 7980
rect 204350 7910 204650 7980
rect 204850 7910 205150 7980
rect 205350 7910 205650 7980
rect 205850 7910 206150 7980
rect 206350 7910 206650 7980
rect 206850 7910 207150 7980
rect 207350 7910 207650 7980
rect 207850 7910 208000 7980
rect 204000 7900 208000 7910
rect 204000 7880 204120 7900
rect 204380 7880 204620 7900
rect 204880 7880 205120 7900
rect 205380 7880 205620 7900
rect 205880 7880 206120 7900
rect 206380 7880 206620 7900
rect 206880 7880 207120 7900
rect 207380 7880 207620 7900
rect 207880 7880 208000 7900
rect 204000 7850 204100 7880
rect 204000 7650 204020 7850
rect 204090 7650 204100 7850
rect 204000 7620 204100 7650
rect 204400 7850 204600 7880
rect 204400 7650 204410 7850
rect 204480 7650 204520 7850
rect 204590 7650 204600 7850
rect 204400 7620 204600 7650
rect 204900 7850 205100 7880
rect 204900 7650 204910 7850
rect 204980 7650 205020 7850
rect 205090 7650 205100 7850
rect 204900 7620 205100 7650
rect 205400 7850 205600 7880
rect 205400 7650 205410 7850
rect 205480 7650 205520 7850
rect 205590 7650 205600 7850
rect 205400 7620 205600 7650
rect 205900 7850 206100 7880
rect 205900 7650 205910 7850
rect 205980 7650 206020 7850
rect 206090 7650 206100 7850
rect 205900 7620 206100 7650
rect 206400 7850 206600 7880
rect 206400 7650 206410 7850
rect 206480 7650 206520 7850
rect 206590 7650 206600 7850
rect 206400 7620 206600 7650
rect 206900 7850 207100 7880
rect 206900 7650 206910 7850
rect 206980 7650 207020 7850
rect 207090 7650 207100 7850
rect 206900 7620 207100 7650
rect 207400 7850 207600 7880
rect 207400 7650 207410 7850
rect 207480 7650 207520 7850
rect 207590 7650 207600 7850
rect 207400 7620 207600 7650
rect 207900 7850 208000 7880
rect 207900 7650 207910 7850
rect 207980 7650 208000 7850
rect 207900 7620 208000 7650
rect 204000 7600 204120 7620
rect 204380 7600 204620 7620
rect 204880 7600 205120 7620
rect 205380 7600 205620 7620
rect 205880 7600 206120 7620
rect 206380 7600 206620 7620
rect 206880 7600 207120 7620
rect 207380 7600 207620 7620
rect 207880 7600 208000 7620
rect 204000 7590 208000 7600
rect 204000 7520 204150 7590
rect 204350 7520 204650 7590
rect 204850 7520 205150 7590
rect 205350 7520 205650 7590
rect 205850 7520 206150 7590
rect 206350 7520 206650 7590
rect 206850 7520 207150 7590
rect 207350 7520 207650 7590
rect 207850 7520 208000 7590
rect 204000 7480 208000 7520
rect 204000 7410 204150 7480
rect 204350 7410 204650 7480
rect 204850 7410 205150 7480
rect 205350 7410 205650 7480
rect 205850 7410 206150 7480
rect 206350 7410 206650 7480
rect 206850 7410 207150 7480
rect 207350 7410 207650 7480
rect 207850 7410 208000 7480
rect 204000 7400 208000 7410
rect 204000 7380 204120 7400
rect 204380 7380 204620 7400
rect 204880 7380 205120 7400
rect 205380 7380 205620 7400
rect 205880 7380 206120 7400
rect 206380 7380 206620 7400
rect 206880 7380 207120 7400
rect 207380 7380 207620 7400
rect 207880 7380 208000 7400
rect 204000 7350 204100 7380
rect 204000 7150 204020 7350
rect 204090 7150 204100 7350
rect 204000 7120 204100 7150
rect 204400 7350 204600 7380
rect 204400 7150 204410 7350
rect 204480 7150 204520 7350
rect 204590 7150 204600 7350
rect 204400 7120 204600 7150
rect 204900 7350 205100 7380
rect 204900 7150 204910 7350
rect 204980 7150 205020 7350
rect 205090 7150 205100 7350
rect 204900 7120 205100 7150
rect 205400 7350 205600 7380
rect 205400 7150 205410 7350
rect 205480 7150 205520 7350
rect 205590 7150 205600 7350
rect 205400 7120 205600 7150
rect 205900 7350 206100 7380
rect 205900 7150 205910 7350
rect 205980 7150 206020 7350
rect 206090 7150 206100 7350
rect 205900 7120 206100 7150
rect 206400 7350 206600 7380
rect 206400 7150 206410 7350
rect 206480 7150 206520 7350
rect 206590 7150 206600 7350
rect 206400 7120 206600 7150
rect 206900 7350 207100 7380
rect 206900 7150 206910 7350
rect 206980 7150 207020 7350
rect 207090 7150 207100 7350
rect 206900 7120 207100 7150
rect 207400 7350 207600 7380
rect 207400 7150 207410 7350
rect 207480 7150 207520 7350
rect 207590 7150 207600 7350
rect 207400 7120 207600 7150
rect 207900 7350 208000 7380
rect 207900 7150 207910 7350
rect 207980 7150 208000 7350
rect 207900 7120 208000 7150
rect 204000 7100 204120 7120
rect 204380 7100 204620 7120
rect 204880 7100 205120 7120
rect 205380 7100 205620 7120
rect 205880 7100 206120 7120
rect 206380 7100 206620 7120
rect 206880 7100 207120 7120
rect 207380 7100 207620 7120
rect 207880 7100 208000 7120
rect 204000 7090 208000 7100
rect 204000 7020 204150 7090
rect 204350 7020 204650 7090
rect 204850 7020 205150 7090
rect 205350 7020 205650 7090
rect 205850 7020 206150 7090
rect 206350 7020 206650 7090
rect 206850 7020 207150 7090
rect 207350 7020 207650 7090
rect 207850 7020 208000 7090
rect 204000 6980 208000 7020
rect 204000 6910 204150 6980
rect 204350 6910 204650 6980
rect 204850 6910 205150 6980
rect 205350 6910 205650 6980
rect 205850 6910 206150 6980
rect 206350 6910 206650 6980
rect 206850 6910 207150 6980
rect 207350 6910 207650 6980
rect 207850 6910 208000 6980
rect 204000 6900 208000 6910
rect 204000 6880 204120 6900
rect 204380 6880 204620 6900
rect 204880 6880 205120 6900
rect 205380 6880 205620 6900
rect 205880 6880 206120 6900
rect 206380 6880 206620 6900
rect 206880 6880 207120 6900
rect 207380 6880 207620 6900
rect 207880 6880 208000 6900
rect 204000 6850 204100 6880
rect 204000 6650 204020 6850
rect 204090 6650 204100 6850
rect 204000 6620 204100 6650
rect 204400 6850 204600 6880
rect 204400 6650 204410 6850
rect 204480 6650 204520 6850
rect 204590 6650 204600 6850
rect 204400 6620 204600 6650
rect 204900 6850 205100 6880
rect 204900 6650 204910 6850
rect 204980 6650 205020 6850
rect 205090 6650 205100 6850
rect 204900 6620 205100 6650
rect 205400 6850 205600 6880
rect 205400 6650 205410 6850
rect 205480 6650 205520 6850
rect 205590 6650 205600 6850
rect 205400 6620 205600 6650
rect 205900 6850 206100 6880
rect 205900 6650 205910 6850
rect 205980 6650 206020 6850
rect 206090 6650 206100 6850
rect 205900 6620 206100 6650
rect 206400 6850 206600 6880
rect 206400 6650 206410 6850
rect 206480 6650 206520 6850
rect 206590 6650 206600 6850
rect 206400 6620 206600 6650
rect 206900 6850 207100 6880
rect 206900 6650 206910 6850
rect 206980 6650 207020 6850
rect 207090 6650 207100 6850
rect 206900 6620 207100 6650
rect 207400 6850 207600 6880
rect 207400 6650 207410 6850
rect 207480 6650 207520 6850
rect 207590 6650 207600 6850
rect 207400 6620 207600 6650
rect 207900 6850 208000 6880
rect 207900 6650 207910 6850
rect 207980 6650 208000 6850
rect 207900 6620 208000 6650
rect 204000 6600 204120 6620
rect 204380 6600 204620 6620
rect 204880 6600 205120 6620
rect 205380 6600 205620 6620
rect 205880 6600 206120 6620
rect 206380 6600 206620 6620
rect 206880 6600 207120 6620
rect 207380 6600 207620 6620
rect 207880 6600 208000 6620
rect 204000 6590 208000 6600
rect 204000 6520 204150 6590
rect 204350 6520 204650 6590
rect 204850 6520 205150 6590
rect 205350 6520 205650 6590
rect 205850 6520 206150 6590
rect 206350 6520 206650 6590
rect 206850 6520 207150 6590
rect 207350 6520 207650 6590
rect 207850 6520 208000 6590
rect 204000 6480 208000 6520
rect 204000 6410 204150 6480
rect 204350 6410 204650 6480
rect 204850 6410 205150 6480
rect 205350 6410 205650 6480
rect 205850 6410 206150 6480
rect 206350 6410 206650 6480
rect 206850 6410 207150 6480
rect 207350 6410 207650 6480
rect 207850 6410 208000 6480
rect 204000 6400 208000 6410
rect 204000 6380 204120 6400
rect 204380 6380 204620 6400
rect 204880 6380 205120 6400
rect 205380 6380 205620 6400
rect 205880 6380 206120 6400
rect 206380 6380 206620 6400
rect 206880 6380 207120 6400
rect 207380 6380 207620 6400
rect 207880 6380 208000 6400
rect 204000 6350 204100 6380
rect 204000 6150 204020 6350
rect 204090 6150 204100 6350
rect 204000 6120 204100 6150
rect 204400 6350 204600 6380
rect 204400 6150 204410 6350
rect 204480 6150 204520 6350
rect 204590 6150 204600 6350
rect 204400 6120 204600 6150
rect 204900 6350 205100 6380
rect 204900 6150 204910 6350
rect 204980 6150 205020 6350
rect 205090 6150 205100 6350
rect 204900 6120 205100 6150
rect 205400 6350 205600 6380
rect 205400 6150 205410 6350
rect 205480 6150 205520 6350
rect 205590 6150 205600 6350
rect 205400 6120 205600 6150
rect 205900 6350 206100 6380
rect 205900 6150 205910 6350
rect 205980 6150 206020 6350
rect 206090 6150 206100 6350
rect 205900 6120 206100 6150
rect 206400 6350 206600 6380
rect 206400 6150 206410 6350
rect 206480 6150 206520 6350
rect 206590 6150 206600 6350
rect 206400 6120 206600 6150
rect 206900 6350 207100 6380
rect 206900 6150 206910 6350
rect 206980 6150 207020 6350
rect 207090 6150 207100 6350
rect 206900 6120 207100 6150
rect 207400 6350 207600 6380
rect 207400 6150 207410 6350
rect 207480 6150 207520 6350
rect 207590 6150 207600 6350
rect 207400 6120 207600 6150
rect 207900 6350 208000 6380
rect 207900 6150 207910 6350
rect 207980 6150 208000 6350
rect 207900 6120 208000 6150
rect 204000 6100 204120 6120
rect 204380 6100 204620 6120
rect 204880 6100 205120 6120
rect 205380 6100 205620 6120
rect 205880 6100 206120 6120
rect 206380 6100 206620 6120
rect 206880 6100 207120 6120
rect 207380 6100 207620 6120
rect 207880 6100 208000 6120
rect 204000 6090 208000 6100
rect 204000 6020 204150 6090
rect 204350 6020 204650 6090
rect 204850 6020 205150 6090
rect 205350 6020 205650 6090
rect 205850 6020 206150 6090
rect 206350 6020 206650 6090
rect 206850 6020 207150 6090
rect 207350 6020 207650 6090
rect 207850 6020 208000 6090
rect 204000 6000 208000 6020
rect 198000 5980 208000 6000
rect 198000 5910 198150 5980
rect 198350 5910 198650 5980
rect 198850 5910 199150 5980
rect 199350 5910 199650 5980
rect 199850 5910 200150 5980
rect 200350 5910 200650 5980
rect 200850 5910 201150 5980
rect 201350 5910 201650 5980
rect 201850 5910 202150 5980
rect 202350 5910 202650 5980
rect 202850 5910 203150 5980
rect 203350 5910 203650 5980
rect 203850 5910 204150 5980
rect 204350 5910 204650 5980
rect 204850 5910 205150 5980
rect 205350 5910 205650 5980
rect 205850 5910 206150 5980
rect 206350 5910 206650 5980
rect 206850 5910 207150 5980
rect 207350 5910 207650 5980
rect 207850 5910 208000 5980
rect 198000 5900 208000 5910
rect 198000 5880 198120 5900
rect 198380 5880 198620 5900
rect 198880 5880 199120 5900
rect 199380 5880 199620 5900
rect 199880 5880 200120 5900
rect 200380 5880 200620 5900
rect 200880 5880 201120 5900
rect 201380 5880 201620 5900
rect 201880 5880 202120 5900
rect 202380 5880 202620 5900
rect 202880 5880 203120 5900
rect 203380 5880 203620 5900
rect 203880 5880 204120 5900
rect 204380 5880 204620 5900
rect 204880 5880 205120 5900
rect 205380 5880 205620 5900
rect 205880 5880 206120 5900
rect 206380 5880 206620 5900
rect 206880 5880 207120 5900
rect 207380 5880 207620 5900
rect 207880 5880 208000 5900
rect 198000 5850 198100 5880
rect 198000 5650 198020 5850
rect 198090 5650 198100 5850
rect 198000 5620 198100 5650
rect 198400 5850 198600 5880
rect 198400 5650 198410 5850
rect 198480 5650 198520 5850
rect 198590 5650 198600 5850
rect 198400 5620 198600 5650
rect 198900 5850 199100 5880
rect 198900 5650 198910 5850
rect 198980 5650 199020 5850
rect 199090 5650 199100 5850
rect 198900 5620 199100 5650
rect 199400 5850 199600 5880
rect 199400 5650 199410 5850
rect 199480 5650 199520 5850
rect 199590 5650 199600 5850
rect 199400 5620 199600 5650
rect 199900 5850 200100 5880
rect 199900 5650 199910 5850
rect 199980 5650 200020 5850
rect 200090 5650 200100 5850
rect 199900 5620 200100 5650
rect 200400 5850 200600 5880
rect 200400 5650 200410 5850
rect 200480 5650 200520 5850
rect 200590 5650 200600 5850
rect 200400 5620 200600 5650
rect 200900 5850 201100 5880
rect 200900 5650 200910 5850
rect 200980 5650 201020 5850
rect 201090 5650 201100 5850
rect 200900 5620 201100 5650
rect 201400 5850 201600 5880
rect 201400 5650 201410 5850
rect 201480 5650 201520 5850
rect 201590 5650 201600 5850
rect 201400 5620 201600 5650
rect 201900 5850 202100 5880
rect 201900 5650 201910 5850
rect 201980 5650 202020 5850
rect 202090 5650 202100 5850
rect 201900 5620 202100 5650
rect 202400 5850 202600 5880
rect 202400 5650 202410 5850
rect 202480 5650 202520 5850
rect 202590 5650 202600 5850
rect 202400 5620 202600 5650
rect 202900 5850 203100 5880
rect 202900 5650 202910 5850
rect 202980 5650 203020 5850
rect 203090 5650 203100 5850
rect 202900 5620 203100 5650
rect 203400 5850 203600 5880
rect 203400 5650 203410 5850
rect 203480 5650 203520 5850
rect 203590 5650 203600 5850
rect 203400 5620 203600 5650
rect 203900 5850 204100 5880
rect 203900 5650 203910 5850
rect 203980 5650 204020 5850
rect 204090 5650 204100 5850
rect 203900 5620 204100 5650
rect 204400 5850 204600 5880
rect 204400 5650 204410 5850
rect 204480 5650 204520 5850
rect 204590 5650 204600 5850
rect 204400 5620 204600 5650
rect 204900 5850 205100 5880
rect 204900 5650 204910 5850
rect 204980 5650 205020 5850
rect 205090 5650 205100 5850
rect 204900 5620 205100 5650
rect 205400 5850 205600 5880
rect 205400 5650 205410 5850
rect 205480 5650 205520 5850
rect 205590 5650 205600 5850
rect 205400 5620 205600 5650
rect 205900 5850 206100 5880
rect 205900 5650 205910 5850
rect 205980 5650 206020 5850
rect 206090 5650 206100 5850
rect 205900 5620 206100 5650
rect 206400 5850 206600 5880
rect 206400 5650 206410 5850
rect 206480 5650 206520 5850
rect 206590 5650 206600 5850
rect 206400 5620 206600 5650
rect 206900 5850 207100 5880
rect 206900 5650 206910 5850
rect 206980 5650 207020 5850
rect 207090 5650 207100 5850
rect 206900 5620 207100 5650
rect 207400 5850 207600 5880
rect 207400 5650 207410 5850
rect 207480 5650 207520 5850
rect 207590 5650 207600 5850
rect 207400 5620 207600 5650
rect 207900 5850 208000 5880
rect 207900 5650 207910 5850
rect 207980 5650 208000 5850
rect 207900 5620 208000 5650
rect 198000 5600 198120 5620
rect 198380 5600 198620 5620
rect 198880 5600 199120 5620
rect 199380 5600 199620 5620
rect 199880 5600 200120 5620
rect 200380 5600 200620 5620
rect 200880 5600 201120 5620
rect 201380 5600 201620 5620
rect 201880 5600 202120 5620
rect 202380 5600 202620 5620
rect 202880 5600 203120 5620
rect 203380 5600 203620 5620
rect 203880 5600 204120 5620
rect 204380 5600 204620 5620
rect 204880 5600 205120 5620
rect 205380 5600 205620 5620
rect 205880 5600 206120 5620
rect 206380 5600 206620 5620
rect 206880 5600 207120 5620
rect 207380 5600 207620 5620
rect 207880 5600 208000 5620
rect 198000 5590 208000 5600
rect 198000 5520 198150 5590
rect 198350 5520 198650 5590
rect 198850 5520 199150 5590
rect 199350 5520 199650 5590
rect 199850 5520 200150 5590
rect 200350 5520 200650 5590
rect 200850 5520 201150 5590
rect 201350 5520 201650 5590
rect 201850 5520 202150 5590
rect 202350 5520 202650 5590
rect 202850 5520 203150 5590
rect 203350 5520 203650 5590
rect 203850 5520 204150 5590
rect 204350 5520 204650 5590
rect 204850 5520 205150 5590
rect 205350 5520 205650 5590
rect 205850 5520 206150 5590
rect 206350 5520 206650 5590
rect 206850 5520 207150 5590
rect 207350 5520 207650 5590
rect 207850 5520 208000 5590
rect 198000 5480 208000 5520
rect 198000 5410 198150 5480
rect 198350 5410 198650 5480
rect 198850 5410 199150 5480
rect 199350 5410 199650 5480
rect 199850 5410 200150 5480
rect 200350 5410 200650 5480
rect 200850 5410 201150 5480
rect 201350 5410 201650 5480
rect 201850 5410 202150 5480
rect 202350 5410 202650 5480
rect 202850 5410 203150 5480
rect 203350 5410 203650 5480
rect 203850 5410 204150 5480
rect 204350 5410 204650 5480
rect 204850 5410 205150 5480
rect 205350 5410 205650 5480
rect 205850 5410 206150 5480
rect 206350 5410 206650 5480
rect 206850 5410 207150 5480
rect 207350 5410 207650 5480
rect 207850 5410 208000 5480
rect 198000 5400 208000 5410
rect 198000 5380 198120 5400
rect 198380 5380 198620 5400
rect 198880 5380 199120 5400
rect 199380 5380 199620 5400
rect 199880 5380 200120 5400
rect 200380 5380 200620 5400
rect 200880 5380 201120 5400
rect 201380 5380 201620 5400
rect 201880 5380 202120 5400
rect 202380 5380 202620 5400
rect 202880 5380 203120 5400
rect 203380 5380 203620 5400
rect 203880 5380 204120 5400
rect 204380 5380 204620 5400
rect 204880 5380 205120 5400
rect 205380 5380 205620 5400
rect 205880 5380 206120 5400
rect 206380 5380 206620 5400
rect 206880 5380 207120 5400
rect 207380 5380 207620 5400
rect 207880 5380 208000 5400
rect 198000 5350 198100 5380
rect 198000 5150 198020 5350
rect 198090 5150 198100 5350
rect 198000 5120 198100 5150
rect 198400 5350 198600 5380
rect 198400 5150 198410 5350
rect 198480 5150 198520 5350
rect 198590 5150 198600 5350
rect 198400 5120 198600 5150
rect 198900 5350 199100 5380
rect 198900 5150 198910 5350
rect 198980 5150 199020 5350
rect 199090 5150 199100 5350
rect 198900 5120 199100 5150
rect 199400 5350 199600 5380
rect 199400 5150 199410 5350
rect 199480 5150 199520 5350
rect 199590 5150 199600 5350
rect 199400 5120 199600 5150
rect 199900 5350 200100 5380
rect 199900 5150 199910 5350
rect 199980 5150 200020 5350
rect 200090 5150 200100 5350
rect 199900 5120 200100 5150
rect 200400 5350 200600 5380
rect 200400 5150 200410 5350
rect 200480 5150 200520 5350
rect 200590 5150 200600 5350
rect 200400 5120 200600 5150
rect 200900 5350 201100 5380
rect 200900 5150 200910 5350
rect 200980 5150 201020 5350
rect 201090 5150 201100 5350
rect 200900 5120 201100 5150
rect 201400 5350 201600 5380
rect 201400 5150 201410 5350
rect 201480 5150 201520 5350
rect 201590 5150 201600 5350
rect 201400 5120 201600 5150
rect 201900 5350 202100 5380
rect 201900 5150 201910 5350
rect 201980 5150 202020 5350
rect 202090 5150 202100 5350
rect 201900 5120 202100 5150
rect 202400 5350 202600 5380
rect 202400 5150 202410 5350
rect 202480 5150 202520 5350
rect 202590 5150 202600 5350
rect 202400 5120 202600 5150
rect 202900 5350 203100 5380
rect 202900 5150 202910 5350
rect 202980 5150 203020 5350
rect 203090 5150 203100 5350
rect 202900 5120 203100 5150
rect 203400 5350 203600 5380
rect 203400 5150 203410 5350
rect 203480 5150 203520 5350
rect 203590 5150 203600 5350
rect 203400 5120 203600 5150
rect 203900 5350 204100 5380
rect 203900 5150 203910 5350
rect 203980 5150 204020 5350
rect 204090 5150 204100 5350
rect 203900 5120 204100 5150
rect 204400 5350 204600 5380
rect 204400 5150 204410 5350
rect 204480 5150 204520 5350
rect 204590 5150 204600 5350
rect 204400 5120 204600 5150
rect 204900 5350 205100 5380
rect 204900 5150 204910 5350
rect 204980 5150 205020 5350
rect 205090 5150 205100 5350
rect 204900 5120 205100 5150
rect 205400 5350 205600 5380
rect 205400 5150 205410 5350
rect 205480 5150 205520 5350
rect 205590 5150 205600 5350
rect 205400 5120 205600 5150
rect 205900 5350 206100 5380
rect 205900 5150 205910 5350
rect 205980 5150 206020 5350
rect 206090 5150 206100 5350
rect 205900 5120 206100 5150
rect 206400 5350 206600 5380
rect 206400 5150 206410 5350
rect 206480 5150 206520 5350
rect 206590 5150 206600 5350
rect 206400 5120 206600 5150
rect 206900 5350 207100 5380
rect 206900 5150 206910 5350
rect 206980 5150 207020 5350
rect 207090 5150 207100 5350
rect 206900 5120 207100 5150
rect 207400 5350 207600 5380
rect 207400 5150 207410 5350
rect 207480 5150 207520 5350
rect 207590 5150 207600 5350
rect 207400 5120 207600 5150
rect 207900 5350 208000 5380
rect 207900 5150 207910 5350
rect 207980 5150 208000 5350
rect 207900 5120 208000 5150
rect 198000 5100 198120 5120
rect 198380 5100 198620 5120
rect 198880 5100 199120 5120
rect 199380 5100 199620 5120
rect 199880 5100 200120 5120
rect 200380 5100 200620 5120
rect 200880 5100 201120 5120
rect 201380 5100 201620 5120
rect 201880 5100 202120 5120
rect 202380 5100 202620 5120
rect 202880 5100 203120 5120
rect 203380 5100 203620 5120
rect 203880 5100 204120 5120
rect 204380 5100 204620 5120
rect 204880 5100 205120 5120
rect 205380 5100 205620 5120
rect 205880 5100 206120 5120
rect 206380 5100 206620 5120
rect 206880 5100 207120 5120
rect 207380 5100 207620 5120
rect 207880 5100 208000 5120
rect 198000 5090 208000 5100
rect 198000 5020 198150 5090
rect 198350 5020 198650 5090
rect 198850 5020 199150 5090
rect 199350 5020 199650 5090
rect 199850 5020 200150 5090
rect 200350 5020 200650 5090
rect 200850 5020 201150 5090
rect 201350 5020 201650 5090
rect 201850 5020 202150 5090
rect 202350 5020 202650 5090
rect 202850 5020 203150 5090
rect 203350 5020 203650 5090
rect 203850 5020 204150 5090
rect 204350 5020 204650 5090
rect 204850 5020 205150 5090
rect 205350 5020 205650 5090
rect 205850 5020 206150 5090
rect 206350 5020 206650 5090
rect 206850 5020 207150 5090
rect 207350 5020 207650 5090
rect 207850 5020 208000 5090
rect 198000 4980 208000 5020
rect 198000 4910 198150 4980
rect 198350 4910 198650 4980
rect 198850 4910 199150 4980
rect 199350 4910 199650 4980
rect 199850 4910 200150 4980
rect 200350 4910 200650 4980
rect 200850 4910 201150 4980
rect 201350 4910 201650 4980
rect 201850 4910 202150 4980
rect 202350 4910 202650 4980
rect 202850 4910 203150 4980
rect 203350 4910 203650 4980
rect 203850 4910 204150 4980
rect 204350 4910 204650 4980
rect 204850 4910 205150 4980
rect 205350 4910 205650 4980
rect 205850 4910 206150 4980
rect 206350 4910 206650 4980
rect 206850 4910 207150 4980
rect 207350 4910 207650 4980
rect 207850 4910 208000 4980
rect 198000 4900 208000 4910
rect 198000 4880 198120 4900
rect 198380 4880 198620 4900
rect 198880 4880 199120 4900
rect 199380 4880 199620 4900
rect 199880 4880 200120 4900
rect 200380 4880 200620 4900
rect 200880 4880 201120 4900
rect 201380 4880 201620 4900
rect 201880 4880 202120 4900
rect 202380 4880 202620 4900
rect 202880 4880 203120 4900
rect 203380 4880 203620 4900
rect 203880 4880 204120 4900
rect 204380 4880 204620 4900
rect 204880 4880 205120 4900
rect 205380 4880 205620 4900
rect 205880 4880 206120 4900
rect 206380 4880 206620 4900
rect 206880 4880 207120 4900
rect 207380 4880 207620 4900
rect 207880 4880 208000 4900
rect 198000 4850 198100 4880
rect 198000 4650 198020 4850
rect 198090 4650 198100 4850
rect 198000 4620 198100 4650
rect 198400 4850 198600 4880
rect 198400 4650 198410 4850
rect 198480 4650 198520 4850
rect 198590 4650 198600 4850
rect 198400 4620 198600 4650
rect 198900 4850 199100 4880
rect 198900 4650 198910 4850
rect 198980 4650 199020 4850
rect 199090 4650 199100 4850
rect 198900 4620 199100 4650
rect 199400 4850 199600 4880
rect 199400 4650 199410 4850
rect 199480 4650 199520 4850
rect 199590 4650 199600 4850
rect 199400 4620 199600 4650
rect 199900 4850 200100 4880
rect 199900 4650 199910 4850
rect 199980 4650 200020 4850
rect 200090 4650 200100 4850
rect 199900 4620 200100 4650
rect 200400 4850 200600 4880
rect 200400 4650 200410 4850
rect 200480 4650 200520 4850
rect 200590 4650 200600 4850
rect 200400 4620 200600 4650
rect 200900 4850 201100 4880
rect 200900 4650 200910 4850
rect 200980 4650 201020 4850
rect 201090 4650 201100 4850
rect 200900 4620 201100 4650
rect 201400 4850 201600 4880
rect 201400 4650 201410 4850
rect 201480 4650 201520 4850
rect 201590 4650 201600 4850
rect 201400 4620 201600 4650
rect 201900 4850 202100 4880
rect 201900 4650 201910 4850
rect 201980 4650 202020 4850
rect 202090 4650 202100 4850
rect 201900 4620 202100 4650
rect 202400 4850 202600 4880
rect 202400 4650 202410 4850
rect 202480 4650 202520 4850
rect 202590 4650 202600 4850
rect 202400 4620 202600 4650
rect 202900 4850 203100 4880
rect 202900 4650 202910 4850
rect 202980 4650 203020 4850
rect 203090 4650 203100 4850
rect 202900 4620 203100 4650
rect 203400 4850 203600 4880
rect 203400 4650 203410 4850
rect 203480 4650 203520 4850
rect 203590 4650 203600 4850
rect 203400 4620 203600 4650
rect 203900 4850 204100 4880
rect 203900 4650 203910 4850
rect 203980 4650 204020 4850
rect 204090 4650 204100 4850
rect 203900 4620 204100 4650
rect 204400 4850 204600 4880
rect 204400 4650 204410 4850
rect 204480 4650 204520 4850
rect 204590 4650 204600 4850
rect 204400 4620 204600 4650
rect 204900 4850 205100 4880
rect 204900 4650 204910 4850
rect 204980 4650 205020 4850
rect 205090 4650 205100 4850
rect 204900 4620 205100 4650
rect 205400 4850 205600 4880
rect 205400 4650 205410 4850
rect 205480 4650 205520 4850
rect 205590 4650 205600 4850
rect 205400 4620 205600 4650
rect 205900 4850 206100 4880
rect 205900 4650 205910 4850
rect 205980 4650 206020 4850
rect 206090 4650 206100 4850
rect 205900 4620 206100 4650
rect 206400 4850 206600 4880
rect 206400 4650 206410 4850
rect 206480 4650 206520 4850
rect 206590 4650 206600 4850
rect 206400 4620 206600 4650
rect 206900 4850 207100 4880
rect 206900 4650 206910 4850
rect 206980 4650 207020 4850
rect 207090 4650 207100 4850
rect 206900 4620 207100 4650
rect 207400 4850 207600 4880
rect 207400 4650 207410 4850
rect 207480 4650 207520 4850
rect 207590 4650 207600 4850
rect 207400 4620 207600 4650
rect 207900 4850 208000 4880
rect 207900 4650 207910 4850
rect 207980 4650 208000 4850
rect 207900 4620 208000 4650
rect 198000 4600 198120 4620
rect 198380 4600 198620 4620
rect 198880 4600 199120 4620
rect 199380 4600 199620 4620
rect 199880 4600 200120 4620
rect 200380 4600 200620 4620
rect 200880 4600 201120 4620
rect 201380 4600 201620 4620
rect 201880 4600 202120 4620
rect 202380 4600 202620 4620
rect 202880 4600 203120 4620
rect 203380 4600 203620 4620
rect 203880 4600 204120 4620
rect 204380 4600 204620 4620
rect 204880 4600 205120 4620
rect 205380 4600 205620 4620
rect 205880 4600 206120 4620
rect 206380 4600 206620 4620
rect 206880 4600 207120 4620
rect 207380 4600 207620 4620
rect 207880 4600 208000 4620
rect 198000 4590 208000 4600
rect 198000 4520 198150 4590
rect 198350 4520 198650 4590
rect 198850 4520 199150 4590
rect 199350 4520 199650 4590
rect 199850 4520 200150 4590
rect 200350 4520 200650 4590
rect 200850 4520 201150 4590
rect 201350 4520 201650 4590
rect 201850 4520 202150 4590
rect 202350 4520 202650 4590
rect 202850 4520 203150 4590
rect 203350 4520 203650 4590
rect 203850 4520 204150 4590
rect 204350 4520 204650 4590
rect 204850 4520 205150 4590
rect 205350 4520 205650 4590
rect 205850 4520 206150 4590
rect 206350 4520 206650 4590
rect 206850 4520 207150 4590
rect 207350 4520 207650 4590
rect 207850 4520 208000 4590
rect 198000 4480 208000 4520
rect 198000 4410 198150 4480
rect 198350 4410 198650 4480
rect 198850 4410 199150 4480
rect 199350 4410 199650 4480
rect 199850 4410 200150 4480
rect 200350 4410 200650 4480
rect 200850 4410 201150 4480
rect 201350 4410 201650 4480
rect 201850 4410 202150 4480
rect 202350 4410 202650 4480
rect 202850 4410 203150 4480
rect 203350 4410 203650 4480
rect 203850 4410 204150 4480
rect 204350 4410 204650 4480
rect 204850 4410 205150 4480
rect 205350 4410 205650 4480
rect 205850 4410 206150 4480
rect 206350 4410 206650 4480
rect 206850 4410 207150 4480
rect 207350 4410 207650 4480
rect 207850 4410 208000 4480
rect 198000 4400 208000 4410
rect 198000 4380 198120 4400
rect 198380 4380 198620 4400
rect 198880 4380 199120 4400
rect 199380 4380 199620 4400
rect 199880 4380 200120 4400
rect 200380 4380 200620 4400
rect 200880 4380 201120 4400
rect 201380 4380 201620 4400
rect 201880 4380 202120 4400
rect 202380 4380 202620 4400
rect 202880 4380 203120 4400
rect 203380 4380 203620 4400
rect 203880 4380 204120 4400
rect 204380 4380 204620 4400
rect 204880 4380 205120 4400
rect 205380 4380 205620 4400
rect 205880 4380 206120 4400
rect 206380 4380 206620 4400
rect 206880 4380 207120 4400
rect 207380 4380 207620 4400
rect 207880 4380 208000 4400
rect 198000 4350 198100 4380
rect 198000 4150 198020 4350
rect 198090 4150 198100 4350
rect 198000 4120 198100 4150
rect 198400 4350 198600 4380
rect 198400 4150 198410 4350
rect 198480 4150 198520 4350
rect 198590 4150 198600 4350
rect 198400 4120 198600 4150
rect 198900 4350 199100 4380
rect 198900 4150 198910 4350
rect 198980 4150 199020 4350
rect 199090 4150 199100 4350
rect 198900 4120 199100 4150
rect 199400 4350 199600 4380
rect 199400 4150 199410 4350
rect 199480 4150 199520 4350
rect 199590 4150 199600 4350
rect 199400 4120 199600 4150
rect 199900 4350 200100 4380
rect 199900 4150 199910 4350
rect 199980 4150 200020 4350
rect 200090 4150 200100 4350
rect 199900 4120 200100 4150
rect 200400 4350 200600 4380
rect 200400 4150 200410 4350
rect 200480 4150 200520 4350
rect 200590 4150 200600 4350
rect 200400 4120 200600 4150
rect 200900 4350 201100 4380
rect 200900 4150 200910 4350
rect 200980 4150 201020 4350
rect 201090 4150 201100 4350
rect 200900 4120 201100 4150
rect 201400 4350 201600 4380
rect 201400 4150 201410 4350
rect 201480 4150 201520 4350
rect 201590 4150 201600 4350
rect 201400 4120 201600 4150
rect 201900 4350 202100 4380
rect 201900 4150 201910 4350
rect 201980 4150 202020 4350
rect 202090 4150 202100 4350
rect 201900 4120 202100 4150
rect 202400 4350 202600 4380
rect 202400 4150 202410 4350
rect 202480 4150 202520 4350
rect 202590 4150 202600 4350
rect 202400 4120 202600 4150
rect 202900 4350 203100 4380
rect 202900 4150 202910 4350
rect 202980 4150 203020 4350
rect 203090 4150 203100 4350
rect 202900 4120 203100 4150
rect 203400 4350 203600 4380
rect 203400 4150 203410 4350
rect 203480 4150 203520 4350
rect 203590 4150 203600 4350
rect 203400 4120 203600 4150
rect 203900 4350 204100 4380
rect 203900 4150 203910 4350
rect 203980 4150 204020 4350
rect 204090 4150 204100 4350
rect 203900 4120 204100 4150
rect 204400 4350 204600 4380
rect 204400 4150 204410 4350
rect 204480 4150 204520 4350
rect 204590 4150 204600 4350
rect 204400 4120 204600 4150
rect 204900 4350 205100 4380
rect 204900 4150 204910 4350
rect 204980 4150 205020 4350
rect 205090 4150 205100 4350
rect 204900 4120 205100 4150
rect 205400 4350 205600 4380
rect 205400 4150 205410 4350
rect 205480 4150 205520 4350
rect 205590 4150 205600 4350
rect 205400 4120 205600 4150
rect 205900 4350 206100 4380
rect 205900 4150 205910 4350
rect 205980 4150 206020 4350
rect 206090 4150 206100 4350
rect 205900 4120 206100 4150
rect 206400 4350 206600 4380
rect 206400 4150 206410 4350
rect 206480 4150 206520 4350
rect 206590 4150 206600 4350
rect 206400 4120 206600 4150
rect 206900 4350 207100 4380
rect 206900 4150 206910 4350
rect 206980 4150 207020 4350
rect 207090 4150 207100 4350
rect 206900 4120 207100 4150
rect 207400 4350 207600 4380
rect 207400 4150 207410 4350
rect 207480 4150 207520 4350
rect 207590 4150 207600 4350
rect 207400 4120 207600 4150
rect 207900 4350 208000 4380
rect 207900 4150 207910 4350
rect 207980 4150 208000 4350
rect 207900 4120 208000 4150
rect 198000 4100 198120 4120
rect 198380 4100 198620 4120
rect 198880 4100 199120 4120
rect 199380 4100 199620 4120
rect 199880 4100 200120 4120
rect 200380 4100 200620 4120
rect 200880 4100 201120 4120
rect 201380 4100 201620 4120
rect 201880 4100 202120 4120
rect 202380 4100 202620 4120
rect 202880 4100 203120 4120
rect 203380 4100 203620 4120
rect 203880 4100 204120 4120
rect 204380 4100 204620 4120
rect 204880 4100 205120 4120
rect 205380 4100 205620 4120
rect 205880 4100 206120 4120
rect 206380 4100 206620 4120
rect 206880 4100 207120 4120
rect 207380 4100 207620 4120
rect 207880 4100 208000 4120
rect 198000 4090 208000 4100
rect 198000 4020 198150 4090
rect 198350 4020 198650 4090
rect 198850 4020 199150 4090
rect 199350 4020 199650 4090
rect 199850 4020 200150 4090
rect 200350 4020 200650 4090
rect 200850 4020 201150 4090
rect 201350 4020 201650 4090
rect 201850 4020 202150 4090
rect 202350 4020 202650 4090
rect 202850 4020 203150 4090
rect 203350 4020 203650 4090
rect 203850 4020 204150 4090
rect 204350 4020 204650 4090
rect 204850 4020 205150 4090
rect 205350 4020 205650 4090
rect 205850 4020 206150 4090
rect 206350 4020 206650 4090
rect 206850 4020 207150 4090
rect 207350 4020 207650 4090
rect 207850 4020 208000 4090
rect 198000 3980 208000 4020
rect 198000 3910 198150 3980
rect 198350 3910 198650 3980
rect 198850 3910 199150 3980
rect 199350 3910 199650 3980
rect 199850 3910 200150 3980
rect 200350 3910 200650 3980
rect 200850 3910 201150 3980
rect 201350 3910 201650 3980
rect 201850 3910 202150 3980
rect 202350 3910 202650 3980
rect 202850 3910 203150 3980
rect 203350 3910 203650 3980
rect 203850 3910 204150 3980
rect 204350 3910 204650 3980
rect 204850 3910 205150 3980
rect 205350 3910 205650 3980
rect 205850 3910 206150 3980
rect 206350 3910 206650 3980
rect 206850 3910 207150 3980
rect 207350 3910 207650 3980
rect 207850 3910 208000 3980
rect 198000 3900 208000 3910
rect 198000 3880 198120 3900
rect 198380 3880 198620 3900
rect 198880 3880 199120 3900
rect 199380 3880 199620 3900
rect 199880 3880 200120 3900
rect 200380 3880 200620 3900
rect 200880 3880 201120 3900
rect 201380 3880 201620 3900
rect 201880 3880 202120 3900
rect 202380 3880 202620 3900
rect 202880 3880 203120 3900
rect 203380 3880 203620 3900
rect 203880 3880 204120 3900
rect 204380 3880 204620 3900
rect 204880 3880 205120 3900
rect 205380 3880 205620 3900
rect 205880 3880 206120 3900
rect 206380 3880 206620 3900
rect 206880 3880 207120 3900
rect 207380 3880 207620 3900
rect 207880 3880 208000 3900
rect 198000 3850 198100 3880
rect 198000 3650 198020 3850
rect 198090 3650 198100 3850
rect 198000 3620 198100 3650
rect 198400 3850 198600 3880
rect 198400 3650 198410 3850
rect 198480 3650 198520 3850
rect 198590 3650 198600 3850
rect 198400 3620 198600 3650
rect 198900 3850 199100 3880
rect 198900 3650 198910 3850
rect 198980 3650 199020 3850
rect 199090 3650 199100 3850
rect 198900 3620 199100 3650
rect 199400 3850 199600 3880
rect 199400 3650 199410 3850
rect 199480 3650 199520 3850
rect 199590 3650 199600 3850
rect 199400 3620 199600 3650
rect 199900 3850 200100 3880
rect 199900 3650 199910 3850
rect 199980 3650 200020 3850
rect 200090 3650 200100 3850
rect 199900 3620 200100 3650
rect 200400 3850 200600 3880
rect 200400 3650 200410 3850
rect 200480 3650 200520 3850
rect 200590 3650 200600 3850
rect 200400 3620 200600 3650
rect 200900 3850 201100 3880
rect 200900 3650 200910 3850
rect 200980 3650 201020 3850
rect 201090 3650 201100 3850
rect 200900 3620 201100 3650
rect 201400 3850 201600 3880
rect 201400 3650 201410 3850
rect 201480 3650 201520 3850
rect 201590 3650 201600 3850
rect 201400 3620 201600 3650
rect 201900 3850 202100 3880
rect 201900 3650 201910 3850
rect 201980 3650 202020 3850
rect 202090 3650 202100 3850
rect 201900 3620 202100 3650
rect 202400 3850 202600 3880
rect 202400 3650 202410 3850
rect 202480 3650 202520 3850
rect 202590 3650 202600 3850
rect 202400 3620 202600 3650
rect 202900 3850 203100 3880
rect 202900 3650 202910 3850
rect 202980 3650 203020 3850
rect 203090 3650 203100 3850
rect 202900 3620 203100 3650
rect 203400 3850 203600 3880
rect 203400 3650 203410 3850
rect 203480 3650 203520 3850
rect 203590 3650 203600 3850
rect 203400 3620 203600 3650
rect 203900 3850 204100 3880
rect 203900 3650 203910 3850
rect 203980 3650 204020 3850
rect 204090 3650 204100 3850
rect 203900 3620 204100 3650
rect 204400 3850 204600 3880
rect 204400 3650 204410 3850
rect 204480 3650 204520 3850
rect 204590 3650 204600 3850
rect 204400 3620 204600 3650
rect 204900 3850 205100 3880
rect 204900 3650 204910 3850
rect 204980 3650 205020 3850
rect 205090 3650 205100 3850
rect 204900 3620 205100 3650
rect 205400 3850 205600 3880
rect 205400 3650 205410 3850
rect 205480 3650 205520 3850
rect 205590 3650 205600 3850
rect 205400 3620 205600 3650
rect 205900 3850 206100 3880
rect 205900 3650 205910 3850
rect 205980 3650 206020 3850
rect 206090 3650 206100 3850
rect 205900 3620 206100 3650
rect 206400 3850 206600 3880
rect 206400 3650 206410 3850
rect 206480 3650 206520 3850
rect 206590 3650 206600 3850
rect 206400 3620 206600 3650
rect 206900 3850 207100 3880
rect 206900 3650 206910 3850
rect 206980 3650 207020 3850
rect 207090 3650 207100 3850
rect 206900 3620 207100 3650
rect 207400 3850 207600 3880
rect 207400 3650 207410 3850
rect 207480 3650 207520 3850
rect 207590 3650 207600 3850
rect 207400 3620 207600 3650
rect 207900 3850 208000 3880
rect 207900 3650 207910 3850
rect 207980 3650 208000 3850
rect 207900 3620 208000 3650
rect 198000 3600 198120 3620
rect 198380 3600 198620 3620
rect 198880 3600 199120 3620
rect 199380 3600 199620 3620
rect 199880 3600 200120 3620
rect 200380 3600 200620 3620
rect 200880 3600 201120 3620
rect 201380 3600 201620 3620
rect 201880 3600 202120 3620
rect 202380 3600 202620 3620
rect 202880 3600 203120 3620
rect 203380 3600 203620 3620
rect 203880 3600 204120 3620
rect 204380 3600 204620 3620
rect 204880 3600 205120 3620
rect 205380 3600 205620 3620
rect 205880 3600 206120 3620
rect 206380 3600 206620 3620
rect 206880 3600 207120 3620
rect 207380 3600 207620 3620
rect 207880 3600 208000 3620
rect 198000 3590 208000 3600
rect 198000 3520 198150 3590
rect 198350 3520 198650 3590
rect 198850 3520 199150 3590
rect 199350 3520 199650 3590
rect 199850 3520 200150 3590
rect 200350 3520 200650 3590
rect 200850 3520 201150 3590
rect 201350 3520 201650 3590
rect 201850 3520 202150 3590
rect 202350 3520 202650 3590
rect 202850 3520 203150 3590
rect 203350 3520 203650 3590
rect 203850 3520 204150 3590
rect 204350 3520 204650 3590
rect 204850 3520 205150 3590
rect 205350 3520 205650 3590
rect 205850 3520 206150 3590
rect 206350 3520 206650 3590
rect 206850 3520 207150 3590
rect 207350 3520 207650 3590
rect 207850 3520 208000 3590
rect 198000 3480 208000 3520
rect 198000 3410 198150 3480
rect 198350 3410 198650 3480
rect 198850 3410 199150 3480
rect 199350 3410 199650 3480
rect 199850 3410 200150 3480
rect 200350 3410 200650 3480
rect 200850 3410 201150 3480
rect 201350 3410 201650 3480
rect 201850 3410 202150 3480
rect 202350 3410 202650 3480
rect 202850 3410 203150 3480
rect 203350 3410 203650 3480
rect 203850 3410 204150 3480
rect 204350 3410 204650 3480
rect 204850 3410 205150 3480
rect 205350 3410 205650 3480
rect 205850 3410 206150 3480
rect 206350 3410 206650 3480
rect 206850 3410 207150 3480
rect 207350 3410 207650 3480
rect 207850 3410 208000 3480
rect 198000 3400 208000 3410
rect 198000 3380 198120 3400
rect 198380 3380 198620 3400
rect 198880 3380 199120 3400
rect 199380 3380 199620 3400
rect 199880 3380 200120 3400
rect 200380 3380 200620 3400
rect 200880 3380 201120 3400
rect 201380 3380 201620 3400
rect 201880 3380 202120 3400
rect 202380 3380 202620 3400
rect 202880 3380 203120 3400
rect 203380 3380 203620 3400
rect 203880 3380 204120 3400
rect 204380 3380 204620 3400
rect 204880 3380 205120 3400
rect 205380 3380 205620 3400
rect 205880 3380 206120 3400
rect 206380 3380 206620 3400
rect 206880 3380 207120 3400
rect 207380 3380 207620 3400
rect 207880 3380 208000 3400
rect 198000 3350 198100 3380
rect 198000 3150 198020 3350
rect 198090 3150 198100 3350
rect 198000 3120 198100 3150
rect 198400 3350 198600 3380
rect 198400 3150 198410 3350
rect 198480 3150 198520 3350
rect 198590 3150 198600 3350
rect 198400 3120 198600 3150
rect 198900 3350 199100 3380
rect 198900 3150 198910 3350
rect 198980 3150 199020 3350
rect 199090 3150 199100 3350
rect 198900 3120 199100 3150
rect 199400 3350 199600 3380
rect 199400 3150 199410 3350
rect 199480 3150 199520 3350
rect 199590 3150 199600 3350
rect 199400 3120 199600 3150
rect 199900 3350 200100 3380
rect 199900 3150 199910 3350
rect 199980 3150 200020 3350
rect 200090 3150 200100 3350
rect 199900 3120 200100 3150
rect 200400 3350 200600 3380
rect 200400 3150 200410 3350
rect 200480 3150 200520 3350
rect 200590 3150 200600 3350
rect 200400 3120 200600 3150
rect 200900 3350 201100 3380
rect 200900 3150 200910 3350
rect 200980 3150 201020 3350
rect 201090 3150 201100 3350
rect 200900 3120 201100 3150
rect 201400 3350 201600 3380
rect 201400 3150 201410 3350
rect 201480 3150 201520 3350
rect 201590 3150 201600 3350
rect 201400 3120 201600 3150
rect 201900 3350 202100 3380
rect 201900 3150 201910 3350
rect 201980 3150 202020 3350
rect 202090 3150 202100 3350
rect 201900 3120 202100 3150
rect 202400 3350 202600 3380
rect 202400 3150 202410 3350
rect 202480 3150 202520 3350
rect 202590 3150 202600 3350
rect 202400 3120 202600 3150
rect 202900 3350 203100 3380
rect 202900 3150 202910 3350
rect 202980 3150 203020 3350
rect 203090 3150 203100 3350
rect 202900 3120 203100 3150
rect 203400 3350 203600 3380
rect 203400 3150 203410 3350
rect 203480 3150 203520 3350
rect 203590 3150 203600 3350
rect 203400 3120 203600 3150
rect 203900 3350 204100 3380
rect 203900 3150 203910 3350
rect 203980 3150 204020 3350
rect 204090 3150 204100 3350
rect 203900 3120 204100 3150
rect 204400 3350 204600 3380
rect 204400 3150 204410 3350
rect 204480 3150 204520 3350
rect 204590 3150 204600 3350
rect 204400 3120 204600 3150
rect 204900 3350 205100 3380
rect 204900 3150 204910 3350
rect 204980 3150 205020 3350
rect 205090 3150 205100 3350
rect 204900 3120 205100 3150
rect 205400 3350 205600 3380
rect 205400 3150 205410 3350
rect 205480 3150 205520 3350
rect 205590 3150 205600 3350
rect 205400 3120 205600 3150
rect 205900 3350 206100 3380
rect 205900 3150 205910 3350
rect 205980 3150 206020 3350
rect 206090 3150 206100 3350
rect 205900 3120 206100 3150
rect 206400 3350 206600 3380
rect 206400 3150 206410 3350
rect 206480 3150 206520 3350
rect 206590 3150 206600 3350
rect 206400 3120 206600 3150
rect 206900 3350 207100 3380
rect 206900 3150 206910 3350
rect 206980 3150 207020 3350
rect 207090 3150 207100 3350
rect 206900 3120 207100 3150
rect 207400 3350 207600 3380
rect 207400 3150 207410 3350
rect 207480 3150 207520 3350
rect 207590 3150 207600 3350
rect 207400 3120 207600 3150
rect 207900 3350 208000 3380
rect 207900 3150 207910 3350
rect 207980 3150 208000 3350
rect 207900 3120 208000 3150
rect 198000 3100 198120 3120
rect 198380 3100 198620 3120
rect 198880 3100 199120 3120
rect 199380 3100 199620 3120
rect 199880 3100 200120 3120
rect 200380 3100 200620 3120
rect 200880 3100 201120 3120
rect 201380 3100 201620 3120
rect 201880 3100 202120 3120
rect 202380 3100 202620 3120
rect 202880 3100 203120 3120
rect 203380 3100 203620 3120
rect 203880 3100 204120 3120
rect 204380 3100 204620 3120
rect 204880 3100 205120 3120
rect 205380 3100 205620 3120
rect 205880 3100 206120 3120
rect 206380 3100 206620 3120
rect 206880 3100 207120 3120
rect 207380 3100 207620 3120
rect 207880 3100 208000 3120
rect 198000 3090 208000 3100
rect 198000 3020 198150 3090
rect 198350 3020 198650 3090
rect 198850 3020 199150 3090
rect 199350 3020 199650 3090
rect 199850 3020 200150 3090
rect 200350 3020 200650 3090
rect 200850 3020 201150 3090
rect 201350 3020 201650 3090
rect 201850 3020 202150 3090
rect 202350 3020 202650 3090
rect 202850 3020 203150 3090
rect 203350 3020 203650 3090
rect 203850 3020 204150 3090
rect 204350 3020 204650 3090
rect 204850 3020 205150 3090
rect 205350 3020 205650 3090
rect 205850 3020 206150 3090
rect 206350 3020 206650 3090
rect 206850 3020 207150 3090
rect 207350 3020 207650 3090
rect 207850 3020 208000 3090
rect 198000 2980 208000 3020
rect 198000 2910 198150 2980
rect 198350 2910 198650 2980
rect 198850 2910 199150 2980
rect 199350 2910 199650 2980
rect 199850 2910 200150 2980
rect 200350 2910 200650 2980
rect 200850 2910 201150 2980
rect 201350 2910 201650 2980
rect 201850 2910 202150 2980
rect 202350 2910 202650 2980
rect 202850 2910 203150 2980
rect 203350 2910 203650 2980
rect 203850 2910 204150 2980
rect 204350 2910 204650 2980
rect 204850 2910 205150 2980
rect 205350 2910 205650 2980
rect 205850 2910 206150 2980
rect 206350 2910 206650 2980
rect 206850 2910 207150 2980
rect 207350 2910 207650 2980
rect 207850 2910 208000 2980
rect 198000 2900 208000 2910
rect 198000 2880 198120 2900
rect 198380 2880 198620 2900
rect 198880 2880 199120 2900
rect 199380 2880 199620 2900
rect 199880 2880 200120 2900
rect 200380 2880 200620 2900
rect 200880 2880 201120 2900
rect 201380 2880 201620 2900
rect 201880 2880 202120 2900
rect 202380 2880 202620 2900
rect 202880 2880 203120 2900
rect 203380 2880 203620 2900
rect 203880 2880 204120 2900
rect 204380 2880 204620 2900
rect 204880 2880 205120 2900
rect 205380 2880 205620 2900
rect 205880 2880 206120 2900
rect 206380 2880 206620 2900
rect 206880 2880 207120 2900
rect 207380 2880 207620 2900
rect 207880 2880 208000 2900
rect 198000 2850 198100 2880
rect 198000 2650 198020 2850
rect 198090 2650 198100 2850
rect 198000 2620 198100 2650
rect 198400 2850 198600 2880
rect 198400 2650 198410 2850
rect 198480 2650 198520 2850
rect 198590 2650 198600 2850
rect 198400 2620 198600 2650
rect 198900 2850 199100 2880
rect 198900 2650 198910 2850
rect 198980 2650 199020 2850
rect 199090 2650 199100 2850
rect 198900 2620 199100 2650
rect 199400 2850 199600 2880
rect 199400 2650 199410 2850
rect 199480 2650 199520 2850
rect 199590 2650 199600 2850
rect 199400 2620 199600 2650
rect 199900 2850 200100 2880
rect 199900 2650 199910 2850
rect 199980 2650 200020 2850
rect 200090 2650 200100 2850
rect 199900 2620 200100 2650
rect 200400 2850 200600 2880
rect 200400 2650 200410 2850
rect 200480 2650 200520 2850
rect 200590 2650 200600 2850
rect 200400 2620 200600 2650
rect 200900 2850 201100 2880
rect 200900 2650 200910 2850
rect 200980 2650 201020 2850
rect 201090 2650 201100 2850
rect 200900 2620 201100 2650
rect 201400 2850 201600 2880
rect 201400 2650 201410 2850
rect 201480 2650 201520 2850
rect 201590 2650 201600 2850
rect 201400 2620 201600 2650
rect 201900 2850 202100 2880
rect 201900 2650 201910 2850
rect 201980 2650 202020 2850
rect 202090 2650 202100 2850
rect 201900 2620 202100 2650
rect 202400 2850 202600 2880
rect 202400 2650 202410 2850
rect 202480 2650 202520 2850
rect 202590 2650 202600 2850
rect 202400 2620 202600 2650
rect 202900 2850 203100 2880
rect 202900 2650 202910 2850
rect 202980 2650 203020 2850
rect 203090 2650 203100 2850
rect 202900 2620 203100 2650
rect 203400 2850 203600 2880
rect 203400 2650 203410 2850
rect 203480 2650 203520 2850
rect 203590 2650 203600 2850
rect 203400 2620 203600 2650
rect 203900 2850 204100 2880
rect 203900 2650 203910 2850
rect 203980 2650 204020 2850
rect 204090 2650 204100 2850
rect 203900 2620 204100 2650
rect 204400 2850 204600 2880
rect 204400 2650 204410 2850
rect 204480 2650 204520 2850
rect 204590 2650 204600 2850
rect 204400 2620 204600 2650
rect 204900 2850 205100 2880
rect 204900 2650 204910 2850
rect 204980 2650 205020 2850
rect 205090 2650 205100 2850
rect 204900 2620 205100 2650
rect 205400 2850 205600 2880
rect 205400 2650 205410 2850
rect 205480 2650 205520 2850
rect 205590 2650 205600 2850
rect 205400 2620 205600 2650
rect 205900 2850 206100 2880
rect 205900 2650 205910 2850
rect 205980 2650 206020 2850
rect 206090 2650 206100 2850
rect 205900 2620 206100 2650
rect 206400 2850 206600 2880
rect 206400 2650 206410 2850
rect 206480 2650 206520 2850
rect 206590 2650 206600 2850
rect 206400 2620 206600 2650
rect 206900 2850 207100 2880
rect 206900 2650 206910 2850
rect 206980 2650 207020 2850
rect 207090 2650 207100 2850
rect 206900 2620 207100 2650
rect 207400 2850 207600 2880
rect 207400 2650 207410 2850
rect 207480 2650 207520 2850
rect 207590 2650 207600 2850
rect 207400 2620 207600 2650
rect 207900 2850 208000 2880
rect 207900 2650 207910 2850
rect 207980 2650 208000 2850
rect 207900 2620 208000 2650
rect 198000 2600 198120 2620
rect 198380 2600 198620 2620
rect 198880 2600 199120 2620
rect 199380 2600 199620 2620
rect 199880 2600 200120 2620
rect 200380 2600 200620 2620
rect 200880 2600 201120 2620
rect 201380 2600 201620 2620
rect 201880 2600 202120 2620
rect 202380 2600 202620 2620
rect 202880 2600 203120 2620
rect 203380 2600 203620 2620
rect 203880 2600 204120 2620
rect 204380 2600 204620 2620
rect 204880 2600 205120 2620
rect 205380 2600 205620 2620
rect 205880 2600 206120 2620
rect 206380 2600 206620 2620
rect 206880 2600 207120 2620
rect 207380 2600 207620 2620
rect 207880 2600 208000 2620
rect 198000 2590 208000 2600
rect 198000 2520 198150 2590
rect 198350 2520 198650 2590
rect 198850 2520 199150 2590
rect 199350 2520 199650 2590
rect 199850 2520 200150 2590
rect 200350 2520 200650 2590
rect 200850 2520 201150 2590
rect 201350 2520 201650 2590
rect 201850 2520 202150 2590
rect 202350 2520 202650 2590
rect 202850 2520 203150 2590
rect 203350 2520 203650 2590
rect 203850 2520 204150 2590
rect 204350 2520 204650 2590
rect 204850 2520 205150 2590
rect 205350 2520 205650 2590
rect 205850 2520 206150 2590
rect 206350 2520 206650 2590
rect 206850 2520 207150 2590
rect 207350 2520 207650 2590
rect 207850 2520 208000 2590
rect 198000 2480 208000 2520
rect 198000 2410 198150 2480
rect 198350 2410 198650 2480
rect 198850 2410 199150 2480
rect 199350 2410 199650 2480
rect 199850 2410 200150 2480
rect 200350 2410 200650 2480
rect 200850 2410 201150 2480
rect 201350 2410 201650 2480
rect 201850 2410 202150 2480
rect 202350 2410 202650 2480
rect 202850 2410 203150 2480
rect 203350 2410 203650 2480
rect 203850 2410 204150 2480
rect 204350 2410 204650 2480
rect 204850 2410 205150 2480
rect 205350 2410 205650 2480
rect 205850 2410 206150 2480
rect 206350 2410 206650 2480
rect 206850 2410 207150 2480
rect 207350 2410 207650 2480
rect 207850 2410 208000 2480
rect 198000 2400 208000 2410
rect 198000 2380 198120 2400
rect 198380 2380 198620 2400
rect 198880 2380 199120 2400
rect 199380 2380 199620 2400
rect 199880 2380 200120 2400
rect 200380 2380 200620 2400
rect 200880 2380 201120 2400
rect 201380 2380 201620 2400
rect 201880 2380 202120 2400
rect 202380 2380 202620 2400
rect 202880 2380 203120 2400
rect 203380 2380 203620 2400
rect 203880 2380 204120 2400
rect 204380 2380 204620 2400
rect 204880 2380 205120 2400
rect 205380 2380 205620 2400
rect 205880 2380 206120 2400
rect 206380 2380 206620 2400
rect 206880 2380 207120 2400
rect 207380 2380 207620 2400
rect 207880 2380 208000 2400
rect 198000 2350 198100 2380
rect 198000 2150 198020 2350
rect 198090 2150 198100 2350
rect 198000 2120 198100 2150
rect 198400 2350 198600 2380
rect 198400 2150 198410 2350
rect 198480 2150 198520 2350
rect 198590 2150 198600 2350
rect 198400 2120 198600 2150
rect 198900 2350 199100 2380
rect 198900 2150 198910 2350
rect 198980 2150 199020 2350
rect 199090 2150 199100 2350
rect 198900 2120 199100 2150
rect 199400 2350 199600 2380
rect 199400 2150 199410 2350
rect 199480 2150 199520 2350
rect 199590 2150 199600 2350
rect 199400 2120 199600 2150
rect 199900 2350 200100 2380
rect 199900 2150 199910 2350
rect 199980 2150 200020 2350
rect 200090 2150 200100 2350
rect 199900 2120 200100 2150
rect 200400 2350 200600 2380
rect 200400 2150 200410 2350
rect 200480 2150 200520 2350
rect 200590 2150 200600 2350
rect 200400 2120 200600 2150
rect 200900 2350 201100 2380
rect 200900 2150 200910 2350
rect 200980 2150 201020 2350
rect 201090 2150 201100 2350
rect 200900 2120 201100 2150
rect 201400 2350 201600 2380
rect 201400 2150 201410 2350
rect 201480 2150 201520 2350
rect 201590 2150 201600 2350
rect 201400 2120 201600 2150
rect 201900 2350 202100 2380
rect 201900 2150 201910 2350
rect 201980 2150 202020 2350
rect 202090 2150 202100 2350
rect 201900 2120 202100 2150
rect 202400 2350 202600 2380
rect 202400 2150 202410 2350
rect 202480 2150 202520 2350
rect 202590 2150 202600 2350
rect 202400 2120 202600 2150
rect 202900 2350 203100 2380
rect 202900 2150 202910 2350
rect 202980 2150 203020 2350
rect 203090 2150 203100 2350
rect 202900 2120 203100 2150
rect 203400 2350 203600 2380
rect 203400 2150 203410 2350
rect 203480 2150 203520 2350
rect 203590 2150 203600 2350
rect 203400 2120 203600 2150
rect 203900 2350 204100 2380
rect 203900 2150 203910 2350
rect 203980 2150 204020 2350
rect 204090 2150 204100 2350
rect 203900 2120 204100 2150
rect 204400 2350 204600 2380
rect 204400 2150 204410 2350
rect 204480 2150 204520 2350
rect 204590 2150 204600 2350
rect 204400 2120 204600 2150
rect 204900 2350 205100 2380
rect 204900 2150 204910 2350
rect 204980 2150 205020 2350
rect 205090 2150 205100 2350
rect 204900 2120 205100 2150
rect 205400 2350 205600 2380
rect 205400 2150 205410 2350
rect 205480 2150 205520 2350
rect 205590 2150 205600 2350
rect 205400 2120 205600 2150
rect 205900 2350 206100 2380
rect 205900 2150 205910 2350
rect 205980 2150 206020 2350
rect 206090 2150 206100 2350
rect 205900 2120 206100 2150
rect 206400 2350 206600 2380
rect 206400 2150 206410 2350
rect 206480 2150 206520 2350
rect 206590 2150 206600 2350
rect 206400 2120 206600 2150
rect 206900 2350 207100 2380
rect 206900 2150 206910 2350
rect 206980 2150 207020 2350
rect 207090 2150 207100 2350
rect 206900 2120 207100 2150
rect 207400 2350 207600 2380
rect 207400 2150 207410 2350
rect 207480 2150 207520 2350
rect 207590 2150 207600 2350
rect 207400 2120 207600 2150
rect 207900 2350 208000 2380
rect 207900 2150 207910 2350
rect 207980 2150 208000 2350
rect 207900 2120 208000 2150
rect 198000 2100 198120 2120
rect 198380 2100 198620 2120
rect 198880 2100 199120 2120
rect 199380 2100 199620 2120
rect 199880 2100 200120 2120
rect 200380 2100 200620 2120
rect 200880 2100 201120 2120
rect 201380 2100 201620 2120
rect 201880 2100 202120 2120
rect 202380 2100 202620 2120
rect 202880 2100 203120 2120
rect 203380 2100 203620 2120
rect 203880 2100 204120 2120
rect 204380 2100 204620 2120
rect 204880 2100 205120 2120
rect 205380 2100 205620 2120
rect 205880 2100 206120 2120
rect 206380 2100 206620 2120
rect 206880 2100 207120 2120
rect 207380 2100 207620 2120
rect 207880 2100 208000 2120
rect 198000 2090 208000 2100
rect 198000 2020 198150 2090
rect 198350 2020 198650 2090
rect 198850 2020 199150 2090
rect 199350 2020 199650 2090
rect 199850 2020 200150 2090
rect 200350 2020 200650 2090
rect 200850 2020 201150 2090
rect 201350 2020 201650 2090
rect 201850 2020 202150 2090
rect 202350 2020 202650 2090
rect 202850 2020 203150 2090
rect 203350 2020 203650 2090
rect 203850 2020 204150 2090
rect 204350 2020 204650 2090
rect 204850 2020 205150 2090
rect 205350 2020 205650 2090
rect 205850 2020 206150 2090
rect 206350 2020 206650 2090
rect 206850 2020 207150 2090
rect 207350 2020 207650 2090
rect 207850 2020 208000 2090
rect 198000 2000 208000 2020
<< via1 >>
rect 250750 136740 250890 136750
rect 250510 135260 250570 135910
rect 250750 134420 250760 136740
rect 250760 134420 250840 136740
rect 250840 134420 250890 136740
rect 250750 134410 250890 134420
rect 171200 119600 181800 121800
rect 222700 119500 231900 121900
rect 196150 103910 196350 103980
rect 196650 103910 196850 103980
rect 197150 103910 197350 103980
rect 197650 103910 197850 103980
rect 198150 103910 198350 103980
rect 198650 103910 198850 103980
rect 199150 103910 199350 103980
rect 199650 103910 199850 103980
rect 200150 103910 200350 103980
rect 200650 103910 200850 103980
rect 201150 103910 201350 103980
rect 201650 103910 201850 103980
rect 202150 103910 202350 103980
rect 202650 103910 202850 103980
rect 203150 103910 203350 103980
rect 203650 103910 203850 103980
rect 204150 103910 204350 103980
rect 204650 103910 204850 103980
rect 205150 103910 205350 103980
rect 205650 103910 205850 103980
rect 206150 103910 206350 103980
rect 206650 103910 206850 103980
rect 207150 103910 207350 103980
rect 207650 103910 207850 103980
rect 196020 103650 196090 103850
rect 196410 103650 196480 103850
rect 196520 103650 196590 103850
rect 196910 103650 196980 103850
rect 197020 103650 197090 103850
rect 197410 103650 197480 103850
rect 197520 103650 197590 103850
rect 197910 103650 197980 103850
rect 198020 103650 198090 103850
rect 198410 103650 198480 103850
rect 198520 103650 198590 103850
rect 198910 103650 198980 103850
rect 199020 103650 199090 103850
rect 199410 103650 199480 103850
rect 199520 103650 199590 103850
rect 199910 103650 199980 103850
rect 200020 103650 200090 103850
rect 200410 103650 200480 103850
rect 200520 103650 200590 103850
rect 200910 103650 200980 103850
rect 201020 103650 201090 103850
rect 201410 103650 201480 103850
rect 201520 103650 201590 103850
rect 201910 103650 201980 103850
rect 202020 103650 202090 103850
rect 202410 103650 202480 103850
rect 202520 103650 202590 103850
rect 202910 103650 202980 103850
rect 203020 103650 203090 103850
rect 203410 103650 203480 103850
rect 203520 103650 203590 103850
rect 203910 103650 203980 103850
rect 204020 103650 204090 103850
rect 204410 103650 204480 103850
rect 204520 103650 204590 103850
rect 204910 103650 204980 103850
rect 205020 103650 205090 103850
rect 205410 103650 205480 103850
rect 205520 103650 205590 103850
rect 205910 103650 205980 103850
rect 206020 103650 206090 103850
rect 206410 103650 206480 103850
rect 206520 103650 206590 103850
rect 206910 103650 206980 103850
rect 207020 103650 207090 103850
rect 207410 103650 207480 103850
rect 207520 103650 207590 103850
rect 207910 103650 207980 103850
rect 196150 103520 196350 103590
rect 196650 103520 196850 103590
rect 197150 103520 197350 103590
rect 197650 103520 197850 103590
rect 198150 103520 198350 103590
rect 198650 103520 198850 103590
rect 199150 103520 199350 103590
rect 199650 103520 199850 103590
rect 200150 103520 200350 103590
rect 200650 103520 200850 103590
rect 201150 103520 201350 103590
rect 201650 103520 201850 103590
rect 202150 103520 202350 103590
rect 202650 103520 202850 103590
rect 203150 103520 203350 103590
rect 203650 103520 203850 103590
rect 204150 103520 204350 103590
rect 204650 103520 204850 103590
rect 205150 103520 205350 103590
rect 205650 103520 205850 103590
rect 206150 103520 206350 103590
rect 206650 103520 206850 103590
rect 207150 103520 207350 103590
rect 207650 103520 207850 103590
rect 196150 103410 196350 103480
rect 196650 103410 196850 103480
rect 197150 103410 197350 103480
rect 197650 103410 197850 103480
rect 198150 103410 198350 103480
rect 198650 103410 198850 103480
rect 199150 103410 199350 103480
rect 199650 103410 199850 103480
rect 200150 103410 200350 103480
rect 200650 103410 200850 103480
rect 201150 103410 201350 103480
rect 201650 103410 201850 103480
rect 202150 103410 202350 103480
rect 202650 103410 202850 103480
rect 203150 103410 203350 103480
rect 203650 103410 203850 103480
rect 204150 103410 204350 103480
rect 204650 103410 204850 103480
rect 205150 103410 205350 103480
rect 205650 103410 205850 103480
rect 206150 103410 206350 103480
rect 206650 103410 206850 103480
rect 207150 103410 207350 103480
rect 207650 103410 207850 103480
rect 196020 103150 196090 103350
rect 196410 103150 196480 103350
rect 196520 103150 196590 103350
rect 196910 103150 196980 103350
rect 197020 103150 197090 103350
rect 197410 103150 197480 103350
rect 197520 103150 197590 103350
rect 197910 103150 197980 103350
rect 198020 103150 198090 103350
rect 198410 103150 198480 103350
rect 198520 103150 198590 103350
rect 198910 103150 198980 103350
rect 199020 103150 199090 103350
rect 199410 103150 199480 103350
rect 199520 103150 199590 103350
rect 199910 103150 199980 103350
rect 200020 103150 200090 103350
rect 200410 103150 200480 103350
rect 200520 103150 200590 103350
rect 200910 103150 200980 103350
rect 201020 103150 201090 103350
rect 201410 103150 201480 103350
rect 201520 103150 201590 103350
rect 201910 103150 201980 103350
rect 202020 103150 202090 103350
rect 202410 103150 202480 103350
rect 202520 103150 202590 103350
rect 202910 103150 202980 103350
rect 203020 103150 203090 103350
rect 203410 103150 203480 103350
rect 203520 103150 203590 103350
rect 203910 103150 203980 103350
rect 204020 103150 204090 103350
rect 204410 103150 204480 103350
rect 204520 103150 204590 103350
rect 204910 103150 204980 103350
rect 205020 103150 205090 103350
rect 205410 103150 205480 103350
rect 205520 103150 205590 103350
rect 205910 103150 205980 103350
rect 206020 103150 206090 103350
rect 206410 103150 206480 103350
rect 206520 103150 206590 103350
rect 206910 103150 206980 103350
rect 207020 103150 207090 103350
rect 207410 103150 207480 103350
rect 207520 103150 207590 103350
rect 207910 103150 207980 103350
rect 196150 103020 196350 103090
rect 196650 103020 196850 103090
rect 197150 103020 197350 103090
rect 197650 103020 197850 103090
rect 198150 103020 198350 103090
rect 198650 103020 198850 103090
rect 199150 103020 199350 103090
rect 199650 103020 199850 103090
rect 200150 103020 200350 103090
rect 200650 103020 200850 103090
rect 201150 103020 201350 103090
rect 201650 103020 201850 103090
rect 202150 103020 202350 103090
rect 202650 103020 202850 103090
rect 203150 103020 203350 103090
rect 203650 103020 203850 103090
rect 204150 103020 204350 103090
rect 204650 103020 204850 103090
rect 205150 103020 205350 103090
rect 205650 103020 205850 103090
rect 206150 103020 206350 103090
rect 206650 103020 206850 103090
rect 207150 103020 207350 103090
rect 207650 103020 207850 103090
rect 196150 102910 196350 102980
rect 196650 102910 196850 102980
rect 197150 102910 197350 102980
rect 197650 102910 197850 102980
rect 198150 102910 198350 102980
rect 198650 102910 198850 102980
rect 199150 102910 199350 102980
rect 199650 102910 199850 102980
rect 200150 102910 200350 102980
rect 200650 102910 200850 102980
rect 201150 102910 201350 102980
rect 201650 102910 201850 102980
rect 202150 102910 202350 102980
rect 202650 102910 202850 102980
rect 203150 102910 203350 102980
rect 203650 102910 203850 102980
rect 204150 102910 204350 102980
rect 204650 102910 204850 102980
rect 205150 102910 205350 102980
rect 205650 102910 205850 102980
rect 206150 102910 206350 102980
rect 206650 102910 206850 102980
rect 207150 102910 207350 102980
rect 207650 102910 207850 102980
rect 196020 102650 196090 102850
rect 196410 102650 196480 102850
rect 196520 102650 196590 102850
rect 196910 102650 196980 102850
rect 197020 102650 197090 102850
rect 197410 102650 197480 102850
rect 197520 102650 197590 102850
rect 197910 102650 197980 102850
rect 198020 102650 198090 102850
rect 198410 102650 198480 102850
rect 198520 102650 198590 102850
rect 198910 102650 198980 102850
rect 199020 102650 199090 102850
rect 199410 102650 199480 102850
rect 199520 102650 199590 102850
rect 199910 102650 199980 102850
rect 200020 102650 200090 102850
rect 200410 102650 200480 102850
rect 200520 102650 200590 102850
rect 200910 102650 200980 102850
rect 201020 102650 201090 102850
rect 201410 102650 201480 102850
rect 201520 102650 201590 102850
rect 201910 102650 201980 102850
rect 202020 102650 202090 102850
rect 202410 102650 202480 102850
rect 202520 102650 202590 102850
rect 202910 102650 202980 102850
rect 203020 102650 203090 102850
rect 203410 102650 203480 102850
rect 203520 102650 203590 102850
rect 203910 102650 203980 102850
rect 204020 102650 204090 102850
rect 204410 102650 204480 102850
rect 204520 102650 204590 102850
rect 204910 102650 204980 102850
rect 205020 102650 205090 102850
rect 205410 102650 205480 102850
rect 205520 102650 205590 102850
rect 205910 102650 205980 102850
rect 206020 102650 206090 102850
rect 206410 102650 206480 102850
rect 206520 102650 206590 102850
rect 206910 102650 206980 102850
rect 207020 102650 207090 102850
rect 207410 102650 207480 102850
rect 207520 102650 207590 102850
rect 207910 102650 207980 102850
rect 196150 102520 196350 102590
rect 196650 102520 196850 102590
rect 197150 102520 197350 102590
rect 197650 102520 197850 102590
rect 198150 102520 198350 102590
rect 198650 102520 198850 102590
rect 199150 102520 199350 102590
rect 199650 102520 199850 102590
rect 200150 102520 200350 102590
rect 200650 102520 200850 102590
rect 201150 102520 201350 102590
rect 201650 102520 201850 102590
rect 202150 102520 202350 102590
rect 202650 102520 202850 102590
rect 203150 102520 203350 102590
rect 203650 102520 203850 102590
rect 204150 102520 204350 102590
rect 204650 102520 204850 102590
rect 205150 102520 205350 102590
rect 205650 102520 205850 102590
rect 206150 102520 206350 102590
rect 206650 102520 206850 102590
rect 207150 102520 207350 102590
rect 207650 102520 207850 102590
rect 196150 102410 196350 102480
rect 196650 102410 196850 102480
rect 197150 102410 197350 102480
rect 197650 102410 197850 102480
rect 198150 102410 198350 102480
rect 198650 102410 198850 102480
rect 199150 102410 199350 102480
rect 199650 102410 199850 102480
rect 200150 102410 200350 102480
rect 200650 102410 200850 102480
rect 201150 102410 201350 102480
rect 201650 102410 201850 102480
rect 202150 102410 202350 102480
rect 202650 102410 202850 102480
rect 203150 102410 203350 102480
rect 203650 102410 203850 102480
rect 204150 102410 204350 102480
rect 204650 102410 204850 102480
rect 205150 102410 205350 102480
rect 205650 102410 205850 102480
rect 206150 102410 206350 102480
rect 206650 102410 206850 102480
rect 207150 102410 207350 102480
rect 207650 102410 207850 102480
rect 196020 102150 196090 102350
rect 196410 102150 196480 102350
rect 196520 102150 196590 102350
rect 196910 102150 196980 102350
rect 197020 102150 197090 102350
rect 197410 102150 197480 102350
rect 197520 102150 197590 102350
rect 197910 102150 197980 102350
rect 198020 102150 198090 102350
rect 198410 102150 198480 102350
rect 198520 102150 198590 102350
rect 198910 102150 198980 102350
rect 199020 102150 199090 102350
rect 199410 102150 199480 102350
rect 199520 102150 199590 102350
rect 199910 102150 199980 102350
rect 200020 102150 200090 102350
rect 200410 102150 200480 102350
rect 200520 102150 200590 102350
rect 200910 102150 200980 102350
rect 201020 102150 201090 102350
rect 201410 102150 201480 102350
rect 201520 102150 201590 102350
rect 201910 102150 201980 102350
rect 202020 102150 202090 102350
rect 202410 102150 202480 102350
rect 202520 102150 202590 102350
rect 202910 102150 202980 102350
rect 203020 102150 203090 102350
rect 203410 102150 203480 102350
rect 203520 102150 203590 102350
rect 203910 102150 203980 102350
rect 204020 102150 204090 102350
rect 204410 102150 204480 102350
rect 204520 102150 204590 102350
rect 204910 102150 204980 102350
rect 205020 102150 205090 102350
rect 205410 102150 205480 102350
rect 205520 102150 205590 102350
rect 205910 102150 205980 102350
rect 206020 102150 206090 102350
rect 206410 102150 206480 102350
rect 206520 102150 206590 102350
rect 206910 102150 206980 102350
rect 207020 102150 207090 102350
rect 207410 102150 207480 102350
rect 207520 102150 207590 102350
rect 207910 102150 207980 102350
rect 196150 102020 196350 102090
rect 196650 102020 196850 102090
rect 197150 102020 197350 102090
rect 197650 102020 197850 102090
rect 198150 102020 198350 102090
rect 198650 102020 198850 102090
rect 199150 102020 199350 102090
rect 199650 102020 199850 102090
rect 200150 102020 200350 102090
rect 200650 102020 200850 102090
rect 201150 102020 201350 102090
rect 201650 102020 201850 102090
rect 202150 102020 202350 102090
rect 202650 102020 202850 102090
rect 203150 102020 203350 102090
rect 203650 102020 203850 102090
rect 204150 102020 204350 102090
rect 204650 102020 204850 102090
rect 205150 102020 205350 102090
rect 205650 102020 205850 102090
rect 206150 102020 206350 102090
rect 206650 102020 206850 102090
rect 207150 102020 207350 102090
rect 207650 102020 207850 102090
rect 196150 101910 196350 101980
rect 196650 101910 196850 101980
rect 197150 101910 197350 101980
rect 197650 101910 197850 101980
rect 198150 101910 198350 101980
rect 198650 101910 198850 101980
rect 199150 101910 199350 101980
rect 199650 101910 199850 101980
rect 200150 101910 200350 101980
rect 200650 101910 200850 101980
rect 201150 101910 201350 101980
rect 201650 101910 201850 101980
rect 202150 101910 202350 101980
rect 202650 101910 202850 101980
rect 203150 101910 203350 101980
rect 203650 101910 203850 101980
rect 204150 101910 204350 101980
rect 204650 101910 204850 101980
rect 205150 101910 205350 101980
rect 205650 101910 205850 101980
rect 206150 101910 206350 101980
rect 206650 101910 206850 101980
rect 207150 101910 207350 101980
rect 207650 101910 207850 101980
rect 196020 101650 196090 101850
rect 196410 101650 196480 101850
rect 196520 101650 196590 101850
rect 196910 101650 196980 101850
rect 197020 101650 197090 101850
rect 197410 101650 197480 101850
rect 197520 101650 197590 101850
rect 197910 101650 197980 101850
rect 198020 101650 198090 101850
rect 198410 101650 198480 101850
rect 198520 101650 198590 101850
rect 198910 101650 198980 101850
rect 199020 101650 199090 101850
rect 199410 101650 199480 101850
rect 199520 101650 199590 101850
rect 199910 101650 199980 101850
rect 200020 101650 200090 101850
rect 200410 101650 200480 101850
rect 200520 101650 200590 101850
rect 200910 101650 200980 101850
rect 201020 101650 201090 101850
rect 201410 101650 201480 101850
rect 201520 101650 201590 101850
rect 201910 101650 201980 101850
rect 202020 101650 202090 101850
rect 202410 101650 202480 101850
rect 202520 101650 202590 101850
rect 202910 101650 202980 101850
rect 203020 101650 203090 101850
rect 203410 101650 203480 101850
rect 203520 101650 203590 101850
rect 203910 101650 203980 101850
rect 204020 101650 204090 101850
rect 204410 101650 204480 101850
rect 204520 101650 204590 101850
rect 204910 101650 204980 101850
rect 205020 101650 205090 101850
rect 205410 101650 205480 101850
rect 205520 101650 205590 101850
rect 205910 101650 205980 101850
rect 206020 101650 206090 101850
rect 206410 101650 206480 101850
rect 206520 101650 206590 101850
rect 206910 101650 206980 101850
rect 207020 101650 207090 101850
rect 207410 101650 207480 101850
rect 207520 101650 207590 101850
rect 207910 101650 207980 101850
rect 196150 101520 196350 101590
rect 196650 101520 196850 101590
rect 197150 101520 197350 101590
rect 197650 101520 197850 101590
rect 198150 101520 198350 101590
rect 198650 101520 198850 101590
rect 199150 101520 199350 101590
rect 199650 101520 199850 101590
rect 200150 101520 200350 101590
rect 200650 101520 200850 101590
rect 201150 101520 201350 101590
rect 201650 101520 201850 101590
rect 202150 101520 202350 101590
rect 202650 101520 202850 101590
rect 203150 101520 203350 101590
rect 203650 101520 203850 101590
rect 204150 101520 204350 101590
rect 204650 101520 204850 101590
rect 205150 101520 205350 101590
rect 205650 101520 205850 101590
rect 206150 101520 206350 101590
rect 206650 101520 206850 101590
rect 207150 101520 207350 101590
rect 207650 101520 207850 101590
rect 196150 101410 196350 101480
rect 196650 101410 196850 101480
rect 197150 101410 197350 101480
rect 197650 101410 197850 101480
rect 198150 101410 198350 101480
rect 198650 101410 198850 101480
rect 199150 101410 199350 101480
rect 199650 101410 199850 101480
rect 200150 101410 200350 101480
rect 200650 101410 200850 101480
rect 201150 101410 201350 101480
rect 201650 101410 201850 101480
rect 202150 101410 202350 101480
rect 202650 101410 202850 101480
rect 203150 101410 203350 101480
rect 203650 101410 203850 101480
rect 204150 101410 204350 101480
rect 204650 101410 204850 101480
rect 205150 101410 205350 101480
rect 205650 101410 205850 101480
rect 206150 101410 206350 101480
rect 206650 101410 206850 101480
rect 207150 101410 207350 101480
rect 207650 101410 207850 101480
rect 196020 101150 196090 101350
rect 196410 101150 196480 101350
rect 196520 101150 196590 101350
rect 196910 101150 196980 101350
rect 197020 101150 197090 101350
rect 197410 101150 197480 101350
rect 197520 101150 197590 101350
rect 197910 101150 197980 101350
rect 198020 101150 198090 101350
rect 198410 101150 198480 101350
rect 198520 101150 198590 101350
rect 198910 101150 198980 101350
rect 199020 101150 199090 101350
rect 199410 101150 199480 101350
rect 199520 101150 199590 101350
rect 199910 101150 199980 101350
rect 200020 101150 200090 101350
rect 200410 101150 200480 101350
rect 200520 101150 200590 101350
rect 200910 101150 200980 101350
rect 201020 101150 201090 101350
rect 201410 101150 201480 101350
rect 201520 101150 201590 101350
rect 201910 101150 201980 101350
rect 202020 101150 202090 101350
rect 202410 101150 202480 101350
rect 202520 101150 202590 101350
rect 202910 101150 202980 101350
rect 203020 101150 203090 101350
rect 203410 101150 203480 101350
rect 203520 101150 203590 101350
rect 203910 101150 203980 101350
rect 204020 101150 204090 101350
rect 204410 101150 204480 101350
rect 204520 101150 204590 101350
rect 204910 101150 204980 101350
rect 205020 101150 205090 101350
rect 205410 101150 205480 101350
rect 205520 101150 205590 101350
rect 205910 101150 205980 101350
rect 206020 101150 206090 101350
rect 206410 101150 206480 101350
rect 206520 101150 206590 101350
rect 206910 101150 206980 101350
rect 207020 101150 207090 101350
rect 207410 101150 207480 101350
rect 207520 101150 207590 101350
rect 207910 101150 207980 101350
rect 196150 101020 196350 101090
rect 196650 101020 196850 101090
rect 197150 101020 197350 101090
rect 197650 101020 197850 101090
rect 198150 101020 198350 101090
rect 198650 101020 198850 101090
rect 199150 101020 199350 101090
rect 199650 101020 199850 101090
rect 200150 101020 200350 101090
rect 200650 101020 200850 101090
rect 201150 101020 201350 101090
rect 201650 101020 201850 101090
rect 202150 101020 202350 101090
rect 202650 101020 202850 101090
rect 203150 101020 203350 101090
rect 203650 101020 203850 101090
rect 204150 101020 204350 101090
rect 204650 101020 204850 101090
rect 205150 101020 205350 101090
rect 205650 101020 205850 101090
rect 206150 101020 206350 101090
rect 206650 101020 206850 101090
rect 207150 101020 207350 101090
rect 207650 101020 207850 101090
rect 196150 100910 196350 100980
rect 196650 100910 196850 100980
rect 197150 100910 197350 100980
rect 197650 100910 197850 100980
rect 198150 100910 198350 100980
rect 198650 100910 198850 100980
rect 199150 100910 199350 100980
rect 199650 100910 199850 100980
rect 200150 100910 200350 100980
rect 200650 100910 200850 100980
rect 201150 100910 201350 100980
rect 201650 100910 201850 100980
rect 202150 100910 202350 100980
rect 202650 100910 202850 100980
rect 203150 100910 203350 100980
rect 203650 100910 203850 100980
rect 204150 100910 204350 100980
rect 204650 100910 204850 100980
rect 205150 100910 205350 100980
rect 205650 100910 205850 100980
rect 206150 100910 206350 100980
rect 206650 100910 206850 100980
rect 207150 100910 207350 100980
rect 207650 100910 207850 100980
rect 196020 100650 196090 100850
rect 196410 100650 196480 100850
rect 196520 100650 196590 100850
rect 196910 100650 196980 100850
rect 197020 100650 197090 100850
rect 197410 100650 197480 100850
rect 197520 100650 197590 100850
rect 197910 100650 197980 100850
rect 198020 100650 198090 100850
rect 198410 100650 198480 100850
rect 198520 100650 198590 100850
rect 198910 100650 198980 100850
rect 199020 100650 199090 100850
rect 199410 100650 199480 100850
rect 199520 100650 199590 100850
rect 199910 100650 199980 100850
rect 200020 100650 200090 100850
rect 200410 100650 200480 100850
rect 200520 100650 200590 100850
rect 200910 100650 200980 100850
rect 201020 100650 201090 100850
rect 201410 100650 201480 100850
rect 201520 100650 201590 100850
rect 201910 100650 201980 100850
rect 202020 100650 202090 100850
rect 202410 100650 202480 100850
rect 202520 100650 202590 100850
rect 202910 100650 202980 100850
rect 203020 100650 203090 100850
rect 203410 100650 203480 100850
rect 203520 100650 203590 100850
rect 203910 100650 203980 100850
rect 204020 100650 204090 100850
rect 204410 100650 204480 100850
rect 204520 100650 204590 100850
rect 204910 100650 204980 100850
rect 205020 100650 205090 100850
rect 205410 100650 205480 100850
rect 205520 100650 205590 100850
rect 205910 100650 205980 100850
rect 206020 100650 206090 100850
rect 206410 100650 206480 100850
rect 206520 100650 206590 100850
rect 206910 100650 206980 100850
rect 207020 100650 207090 100850
rect 207410 100650 207480 100850
rect 207520 100650 207590 100850
rect 207910 100650 207980 100850
rect 196150 100520 196350 100590
rect 196650 100520 196850 100590
rect 197150 100520 197350 100590
rect 197650 100520 197850 100590
rect 198150 100520 198350 100590
rect 198650 100520 198850 100590
rect 199150 100520 199350 100590
rect 199650 100520 199850 100590
rect 200150 100520 200350 100590
rect 200650 100520 200850 100590
rect 201150 100520 201350 100590
rect 201650 100520 201850 100590
rect 202150 100520 202350 100590
rect 202650 100520 202850 100590
rect 203150 100520 203350 100590
rect 203650 100520 203850 100590
rect 204150 100520 204350 100590
rect 204650 100520 204850 100590
rect 205150 100520 205350 100590
rect 205650 100520 205850 100590
rect 206150 100520 206350 100590
rect 206650 100520 206850 100590
rect 207150 100520 207350 100590
rect 207650 100520 207850 100590
rect 196150 100410 196350 100480
rect 196650 100410 196850 100480
rect 197150 100410 197350 100480
rect 197650 100410 197850 100480
rect 198150 100410 198350 100480
rect 198650 100410 198850 100480
rect 199150 100410 199350 100480
rect 199650 100410 199850 100480
rect 200150 100410 200350 100480
rect 200650 100410 200850 100480
rect 201150 100410 201350 100480
rect 201650 100410 201850 100480
rect 202150 100410 202350 100480
rect 202650 100410 202850 100480
rect 203150 100410 203350 100480
rect 203650 100410 203850 100480
rect 204150 100410 204350 100480
rect 204650 100410 204850 100480
rect 205150 100410 205350 100480
rect 205650 100410 205850 100480
rect 206150 100410 206350 100480
rect 206650 100410 206850 100480
rect 207150 100410 207350 100480
rect 207650 100410 207850 100480
rect 196020 100150 196090 100350
rect 196410 100150 196480 100350
rect 196520 100150 196590 100350
rect 196910 100150 196980 100350
rect 197020 100150 197090 100350
rect 197410 100150 197480 100350
rect 197520 100150 197590 100350
rect 197910 100150 197980 100350
rect 198020 100150 198090 100350
rect 198410 100150 198480 100350
rect 198520 100150 198590 100350
rect 198910 100150 198980 100350
rect 199020 100150 199090 100350
rect 199410 100150 199480 100350
rect 199520 100150 199590 100350
rect 199910 100150 199980 100350
rect 200020 100150 200090 100350
rect 200410 100150 200480 100350
rect 200520 100150 200590 100350
rect 200910 100150 200980 100350
rect 201020 100150 201090 100350
rect 201410 100150 201480 100350
rect 201520 100150 201590 100350
rect 201910 100150 201980 100350
rect 202020 100150 202090 100350
rect 202410 100150 202480 100350
rect 202520 100150 202590 100350
rect 202910 100150 202980 100350
rect 203020 100150 203090 100350
rect 203410 100150 203480 100350
rect 203520 100150 203590 100350
rect 203910 100150 203980 100350
rect 204020 100150 204090 100350
rect 204410 100150 204480 100350
rect 204520 100150 204590 100350
rect 204910 100150 204980 100350
rect 205020 100150 205090 100350
rect 205410 100150 205480 100350
rect 205520 100150 205590 100350
rect 205910 100150 205980 100350
rect 206020 100150 206090 100350
rect 206410 100150 206480 100350
rect 206520 100150 206590 100350
rect 206910 100150 206980 100350
rect 207020 100150 207090 100350
rect 207410 100150 207480 100350
rect 207520 100150 207590 100350
rect 207910 100150 207980 100350
rect 196150 100020 196350 100090
rect 196650 100020 196850 100090
rect 197150 100020 197350 100090
rect 197650 100020 197850 100090
rect 198150 100020 198350 100090
rect 198650 100020 198850 100090
rect 199150 100020 199350 100090
rect 199650 100020 199850 100090
rect 200150 100020 200350 100090
rect 200650 100020 200850 100090
rect 201150 100020 201350 100090
rect 201650 100020 201850 100090
rect 202150 100020 202350 100090
rect 202650 100020 202850 100090
rect 203150 100020 203350 100090
rect 203650 100020 203850 100090
rect 204150 100020 204350 100090
rect 204650 100020 204850 100090
rect 205150 100020 205350 100090
rect 205650 100020 205850 100090
rect 206150 100020 206350 100090
rect 206650 100020 206850 100090
rect 207150 100020 207350 100090
rect 207650 100020 207850 100090
rect 196150 99910 196350 99980
rect 196650 99910 196850 99980
rect 197150 99910 197350 99980
rect 197650 99910 197850 99980
rect 198150 99910 198350 99980
rect 198650 99910 198850 99980
rect 199150 99910 199350 99980
rect 199650 99910 199850 99980
rect 200150 99910 200350 99980
rect 200650 99910 200850 99980
rect 201150 99910 201350 99980
rect 201650 99910 201850 99980
rect 202150 99910 202350 99980
rect 202650 99910 202850 99980
rect 203150 99910 203350 99980
rect 203650 99910 203850 99980
rect 204150 99910 204350 99980
rect 204650 99910 204850 99980
rect 205150 99910 205350 99980
rect 205650 99910 205850 99980
rect 206150 99910 206350 99980
rect 206650 99910 206850 99980
rect 207150 99910 207350 99980
rect 207650 99910 207850 99980
rect 196020 99650 196090 99850
rect 196410 99650 196480 99850
rect 196520 99650 196590 99850
rect 196910 99650 196980 99850
rect 197020 99650 197090 99850
rect 197410 99650 197480 99850
rect 197520 99650 197590 99850
rect 197910 99650 197980 99850
rect 198020 99650 198090 99850
rect 198410 99650 198480 99850
rect 198520 99650 198590 99850
rect 198910 99650 198980 99850
rect 199020 99650 199090 99850
rect 199410 99650 199480 99850
rect 199520 99650 199590 99850
rect 199910 99650 199980 99850
rect 200020 99650 200090 99850
rect 200410 99650 200480 99850
rect 200520 99650 200590 99850
rect 200910 99650 200980 99850
rect 201020 99650 201090 99850
rect 201410 99650 201480 99850
rect 201520 99650 201590 99850
rect 201910 99650 201980 99850
rect 202020 99650 202090 99850
rect 202410 99650 202480 99850
rect 202520 99650 202590 99850
rect 202910 99650 202980 99850
rect 203020 99650 203090 99850
rect 203410 99650 203480 99850
rect 203520 99650 203590 99850
rect 203910 99650 203980 99850
rect 204020 99650 204090 99850
rect 204410 99650 204480 99850
rect 204520 99650 204590 99850
rect 204910 99650 204980 99850
rect 205020 99650 205090 99850
rect 205410 99650 205480 99850
rect 205520 99650 205590 99850
rect 205910 99650 205980 99850
rect 206020 99650 206090 99850
rect 206410 99650 206480 99850
rect 206520 99650 206590 99850
rect 206910 99650 206980 99850
rect 207020 99650 207090 99850
rect 207410 99650 207480 99850
rect 207520 99650 207590 99850
rect 207910 99650 207980 99850
rect 196150 99520 196350 99590
rect 196650 99520 196850 99590
rect 197150 99520 197350 99590
rect 197650 99520 197850 99590
rect 198150 99520 198350 99590
rect 198650 99520 198850 99590
rect 199150 99520 199350 99590
rect 199650 99520 199850 99590
rect 200150 99520 200350 99590
rect 200650 99520 200850 99590
rect 201150 99520 201350 99590
rect 201650 99520 201850 99590
rect 202150 99520 202350 99590
rect 202650 99520 202850 99590
rect 203150 99520 203350 99590
rect 203650 99520 203850 99590
rect 204150 99520 204350 99590
rect 204650 99520 204850 99590
rect 205150 99520 205350 99590
rect 205650 99520 205850 99590
rect 206150 99520 206350 99590
rect 206650 99520 206850 99590
rect 207150 99520 207350 99590
rect 207650 99520 207850 99590
rect 196150 99410 196350 99480
rect 196650 99410 196850 99480
rect 197150 99410 197350 99480
rect 197650 99410 197850 99480
rect 198150 99410 198350 99480
rect 198650 99410 198850 99480
rect 199150 99410 199350 99480
rect 199650 99410 199850 99480
rect 200150 99410 200350 99480
rect 200650 99410 200850 99480
rect 201150 99410 201350 99480
rect 201650 99410 201850 99480
rect 202150 99410 202350 99480
rect 202650 99410 202850 99480
rect 203150 99410 203350 99480
rect 203650 99410 203850 99480
rect 204150 99410 204350 99480
rect 204650 99410 204850 99480
rect 205150 99410 205350 99480
rect 205650 99410 205850 99480
rect 206150 99410 206350 99480
rect 206650 99410 206850 99480
rect 207150 99410 207350 99480
rect 207650 99410 207850 99480
rect 196020 99150 196090 99350
rect 196410 99150 196480 99350
rect 196520 99150 196590 99350
rect 196910 99150 196980 99350
rect 197020 99150 197090 99350
rect 197410 99150 197480 99350
rect 197520 99150 197590 99350
rect 197910 99150 197980 99350
rect 198020 99150 198090 99350
rect 198410 99150 198480 99350
rect 198520 99150 198590 99350
rect 198910 99150 198980 99350
rect 199020 99150 199090 99350
rect 199410 99150 199480 99350
rect 199520 99150 199590 99350
rect 199910 99150 199980 99350
rect 200020 99150 200090 99350
rect 200410 99150 200480 99350
rect 200520 99150 200590 99350
rect 200910 99150 200980 99350
rect 201020 99150 201090 99350
rect 201410 99150 201480 99350
rect 201520 99150 201590 99350
rect 201910 99150 201980 99350
rect 202020 99150 202090 99350
rect 202410 99150 202480 99350
rect 202520 99150 202590 99350
rect 202910 99150 202980 99350
rect 203020 99150 203090 99350
rect 203410 99150 203480 99350
rect 203520 99150 203590 99350
rect 203910 99150 203980 99350
rect 204020 99150 204090 99350
rect 204410 99150 204480 99350
rect 204520 99150 204590 99350
rect 204910 99150 204980 99350
rect 205020 99150 205090 99350
rect 205410 99150 205480 99350
rect 205520 99150 205590 99350
rect 205910 99150 205980 99350
rect 206020 99150 206090 99350
rect 206410 99150 206480 99350
rect 206520 99150 206590 99350
rect 206910 99150 206980 99350
rect 207020 99150 207090 99350
rect 207410 99150 207480 99350
rect 207520 99150 207590 99350
rect 207910 99150 207980 99350
rect 196150 99020 196350 99090
rect 196650 99020 196850 99090
rect 197150 99020 197350 99090
rect 197650 99020 197850 99090
rect 198150 99020 198350 99090
rect 198650 99020 198850 99090
rect 199150 99020 199350 99090
rect 199650 99020 199850 99090
rect 200150 99020 200350 99090
rect 200650 99020 200850 99090
rect 201150 99020 201350 99090
rect 201650 99020 201850 99090
rect 202150 99020 202350 99090
rect 202650 99020 202850 99090
rect 203150 99020 203350 99090
rect 203650 99020 203850 99090
rect 204150 99020 204350 99090
rect 204650 99020 204850 99090
rect 205150 99020 205350 99090
rect 205650 99020 205850 99090
rect 206150 99020 206350 99090
rect 206650 99020 206850 99090
rect 207150 99020 207350 99090
rect 207650 99020 207850 99090
rect 196150 98910 196350 98980
rect 196650 98910 196850 98980
rect 197150 98910 197350 98980
rect 197650 98910 197850 98980
rect 198150 98910 198350 98980
rect 198650 98910 198850 98980
rect 199150 98910 199350 98980
rect 199650 98910 199850 98980
rect 200150 98910 200350 98980
rect 200650 98910 200850 98980
rect 201150 98910 201350 98980
rect 201650 98910 201850 98980
rect 202150 98910 202350 98980
rect 202650 98910 202850 98980
rect 203150 98910 203350 98980
rect 203650 98910 203850 98980
rect 204150 98910 204350 98980
rect 204650 98910 204850 98980
rect 205150 98910 205350 98980
rect 205650 98910 205850 98980
rect 206150 98910 206350 98980
rect 206650 98910 206850 98980
rect 207150 98910 207350 98980
rect 207650 98910 207850 98980
rect 196020 98650 196090 98850
rect 196410 98650 196480 98850
rect 196520 98650 196590 98850
rect 196910 98650 196980 98850
rect 197020 98650 197090 98850
rect 197410 98650 197480 98850
rect 197520 98650 197590 98850
rect 197910 98650 197980 98850
rect 198020 98650 198090 98850
rect 198410 98650 198480 98850
rect 198520 98650 198590 98850
rect 198910 98650 198980 98850
rect 199020 98650 199090 98850
rect 199410 98650 199480 98850
rect 199520 98650 199590 98850
rect 199910 98650 199980 98850
rect 200020 98650 200090 98850
rect 200410 98650 200480 98850
rect 200520 98650 200590 98850
rect 200910 98650 200980 98850
rect 201020 98650 201090 98850
rect 201410 98650 201480 98850
rect 201520 98650 201590 98850
rect 201910 98650 201980 98850
rect 202020 98650 202090 98850
rect 202410 98650 202480 98850
rect 202520 98650 202590 98850
rect 202910 98650 202980 98850
rect 203020 98650 203090 98850
rect 203410 98650 203480 98850
rect 203520 98650 203590 98850
rect 203910 98650 203980 98850
rect 204020 98650 204090 98850
rect 204410 98650 204480 98850
rect 204520 98650 204590 98850
rect 204910 98650 204980 98850
rect 205020 98650 205090 98850
rect 205410 98650 205480 98850
rect 205520 98650 205590 98850
rect 205910 98650 205980 98850
rect 206020 98650 206090 98850
rect 206410 98650 206480 98850
rect 206520 98650 206590 98850
rect 206910 98650 206980 98850
rect 207020 98650 207090 98850
rect 207410 98650 207480 98850
rect 207520 98650 207590 98850
rect 207910 98650 207980 98850
rect 196150 98520 196350 98590
rect 196650 98520 196850 98590
rect 197150 98520 197350 98590
rect 197650 98520 197850 98590
rect 198150 98520 198350 98590
rect 198650 98520 198850 98590
rect 199150 98520 199350 98590
rect 199650 98520 199850 98590
rect 200150 98520 200350 98590
rect 200650 98520 200850 98590
rect 201150 98520 201350 98590
rect 201650 98520 201850 98590
rect 202150 98520 202350 98590
rect 202650 98520 202850 98590
rect 203150 98520 203350 98590
rect 203650 98520 203850 98590
rect 204150 98520 204350 98590
rect 204650 98520 204850 98590
rect 205150 98520 205350 98590
rect 205650 98520 205850 98590
rect 206150 98520 206350 98590
rect 206650 98520 206850 98590
rect 207150 98520 207350 98590
rect 207650 98520 207850 98590
rect 196150 98410 196350 98480
rect 196650 98410 196850 98480
rect 197150 98410 197350 98480
rect 197650 98410 197850 98480
rect 198150 98410 198350 98480
rect 198650 98410 198850 98480
rect 199150 98410 199350 98480
rect 199650 98410 199850 98480
rect 200150 98410 200350 98480
rect 200650 98410 200850 98480
rect 201150 98410 201350 98480
rect 201650 98410 201850 98480
rect 202150 98410 202350 98480
rect 202650 98410 202850 98480
rect 203150 98410 203350 98480
rect 203650 98410 203850 98480
rect 204150 98410 204350 98480
rect 204650 98410 204850 98480
rect 205150 98410 205350 98480
rect 205650 98410 205850 98480
rect 206150 98410 206350 98480
rect 206650 98410 206850 98480
rect 207150 98410 207350 98480
rect 207650 98410 207850 98480
rect 196020 98150 196090 98350
rect 196410 98150 196480 98350
rect 196520 98150 196590 98350
rect 196910 98150 196980 98350
rect 197020 98150 197090 98350
rect 197410 98150 197480 98350
rect 197520 98150 197590 98350
rect 197910 98150 197980 98350
rect 198020 98150 198090 98350
rect 198410 98150 198480 98350
rect 198520 98150 198590 98350
rect 198910 98150 198980 98350
rect 199020 98150 199090 98350
rect 199410 98150 199480 98350
rect 199520 98150 199590 98350
rect 199910 98150 199980 98350
rect 200020 98150 200090 98350
rect 200410 98150 200480 98350
rect 200520 98150 200590 98350
rect 200910 98150 200980 98350
rect 201020 98150 201090 98350
rect 201410 98150 201480 98350
rect 201520 98150 201590 98350
rect 201910 98150 201980 98350
rect 202020 98150 202090 98350
rect 202410 98150 202480 98350
rect 202520 98150 202590 98350
rect 202910 98150 202980 98350
rect 203020 98150 203090 98350
rect 203410 98150 203480 98350
rect 203520 98150 203590 98350
rect 203910 98150 203980 98350
rect 204020 98150 204090 98350
rect 204410 98150 204480 98350
rect 204520 98150 204590 98350
rect 204910 98150 204980 98350
rect 205020 98150 205090 98350
rect 205410 98150 205480 98350
rect 205520 98150 205590 98350
rect 205910 98150 205980 98350
rect 206020 98150 206090 98350
rect 206410 98150 206480 98350
rect 206520 98150 206590 98350
rect 206910 98150 206980 98350
rect 207020 98150 207090 98350
rect 207410 98150 207480 98350
rect 207520 98150 207590 98350
rect 207910 98150 207980 98350
rect 196150 98020 196350 98090
rect 196650 98020 196850 98090
rect 197150 98020 197350 98090
rect 197650 98020 197850 98090
rect 198150 98020 198350 98090
rect 198650 98020 198850 98090
rect 199150 98020 199350 98090
rect 199650 98020 199850 98090
rect 200150 98020 200350 98090
rect 200650 98020 200850 98090
rect 201150 98020 201350 98090
rect 201650 98020 201850 98090
rect 202150 98020 202350 98090
rect 202650 98020 202850 98090
rect 203150 98020 203350 98090
rect 203650 98020 203850 98090
rect 204150 98020 204350 98090
rect 204650 98020 204850 98090
rect 205150 98020 205350 98090
rect 205650 98020 205850 98090
rect 206150 98020 206350 98090
rect 206650 98020 206850 98090
rect 207150 98020 207350 98090
rect 207650 98020 207850 98090
rect 196150 97910 196350 97980
rect 196650 97910 196850 97980
rect 197150 97910 197350 97980
rect 197650 97910 197850 97980
rect 198150 97910 198350 97980
rect 198650 97910 198850 97980
rect 199150 97910 199350 97980
rect 199650 97910 199850 97980
rect 200150 97910 200350 97980
rect 200650 97910 200850 97980
rect 201150 97910 201350 97980
rect 201650 97910 201850 97980
rect 202150 97910 202350 97980
rect 202650 97910 202850 97980
rect 203150 97910 203350 97980
rect 203650 97910 203850 97980
rect 204150 97910 204350 97980
rect 204650 97910 204850 97980
rect 205150 97910 205350 97980
rect 205650 97910 205850 97980
rect 206150 97910 206350 97980
rect 206650 97910 206850 97980
rect 207150 97910 207350 97980
rect 207650 97910 207850 97980
rect 196020 97650 196090 97850
rect 196410 97650 196480 97850
rect 196520 97650 196590 97850
rect 196910 97650 196980 97850
rect 197020 97650 197090 97850
rect 197410 97650 197480 97850
rect 197520 97650 197590 97850
rect 197910 97650 197980 97850
rect 198020 97650 198090 97850
rect 198410 97650 198480 97850
rect 198520 97650 198590 97850
rect 198910 97650 198980 97850
rect 199020 97650 199090 97850
rect 199410 97650 199480 97850
rect 199520 97650 199590 97850
rect 199910 97650 199980 97850
rect 200020 97650 200090 97850
rect 200410 97650 200480 97850
rect 200520 97650 200590 97850
rect 200910 97650 200980 97850
rect 201020 97650 201090 97850
rect 201410 97650 201480 97850
rect 201520 97650 201590 97850
rect 201910 97650 201980 97850
rect 202020 97650 202090 97850
rect 202410 97650 202480 97850
rect 202520 97650 202590 97850
rect 202910 97650 202980 97850
rect 203020 97650 203090 97850
rect 203410 97650 203480 97850
rect 203520 97650 203590 97850
rect 203910 97650 203980 97850
rect 204020 97650 204090 97850
rect 204410 97650 204480 97850
rect 204520 97650 204590 97850
rect 204910 97650 204980 97850
rect 205020 97650 205090 97850
rect 205410 97650 205480 97850
rect 205520 97650 205590 97850
rect 205910 97650 205980 97850
rect 206020 97650 206090 97850
rect 206410 97650 206480 97850
rect 206520 97650 206590 97850
rect 206910 97650 206980 97850
rect 207020 97650 207090 97850
rect 207410 97650 207480 97850
rect 207520 97650 207590 97850
rect 207910 97650 207980 97850
rect 196150 97520 196350 97590
rect 196650 97520 196850 97590
rect 197150 97520 197350 97590
rect 197650 97520 197850 97590
rect 198150 97520 198350 97590
rect 198650 97520 198850 97590
rect 199150 97520 199350 97590
rect 199650 97520 199850 97590
rect 200150 97520 200350 97590
rect 200650 97520 200850 97590
rect 201150 97520 201350 97590
rect 201650 97520 201850 97590
rect 202150 97520 202350 97590
rect 202650 97520 202850 97590
rect 203150 97520 203350 97590
rect 203650 97520 203850 97590
rect 204150 97520 204350 97590
rect 204650 97520 204850 97590
rect 205150 97520 205350 97590
rect 205650 97520 205850 97590
rect 206150 97520 206350 97590
rect 206650 97520 206850 97590
rect 207150 97520 207350 97590
rect 207650 97520 207850 97590
rect 196150 97410 196350 97480
rect 196650 97410 196850 97480
rect 197150 97410 197350 97480
rect 197650 97410 197850 97480
rect 198150 97410 198350 97480
rect 198650 97410 198850 97480
rect 199150 97410 199350 97480
rect 199650 97410 199850 97480
rect 200150 97410 200350 97480
rect 200650 97410 200850 97480
rect 201150 97410 201350 97480
rect 201650 97410 201850 97480
rect 202150 97410 202350 97480
rect 202650 97410 202850 97480
rect 203150 97410 203350 97480
rect 203650 97410 203850 97480
rect 204150 97410 204350 97480
rect 204650 97410 204850 97480
rect 205150 97410 205350 97480
rect 205650 97410 205850 97480
rect 206150 97410 206350 97480
rect 206650 97410 206850 97480
rect 207150 97410 207350 97480
rect 207650 97410 207850 97480
rect 196020 97150 196090 97350
rect 196410 97150 196480 97350
rect 196520 97150 196590 97350
rect 196910 97150 196980 97350
rect 197020 97150 197090 97350
rect 197410 97150 197480 97350
rect 197520 97150 197590 97350
rect 197910 97150 197980 97350
rect 198020 97150 198090 97350
rect 198410 97150 198480 97350
rect 198520 97150 198590 97350
rect 198910 97150 198980 97350
rect 199020 97150 199090 97350
rect 199410 97150 199480 97350
rect 199520 97150 199590 97350
rect 199910 97150 199980 97350
rect 200020 97150 200090 97350
rect 200410 97150 200480 97350
rect 200520 97150 200590 97350
rect 200910 97150 200980 97350
rect 201020 97150 201090 97350
rect 201410 97150 201480 97350
rect 201520 97150 201590 97350
rect 201910 97150 201980 97350
rect 202020 97150 202090 97350
rect 202410 97150 202480 97350
rect 202520 97150 202590 97350
rect 202910 97150 202980 97350
rect 203020 97150 203090 97350
rect 203410 97150 203480 97350
rect 203520 97150 203590 97350
rect 203910 97150 203980 97350
rect 204020 97150 204090 97350
rect 204410 97150 204480 97350
rect 204520 97150 204590 97350
rect 204910 97150 204980 97350
rect 205020 97150 205090 97350
rect 205410 97150 205480 97350
rect 205520 97150 205590 97350
rect 205910 97150 205980 97350
rect 206020 97150 206090 97350
rect 206410 97150 206480 97350
rect 206520 97150 206590 97350
rect 206910 97150 206980 97350
rect 207020 97150 207090 97350
rect 207410 97150 207480 97350
rect 207520 97150 207590 97350
rect 207910 97150 207980 97350
rect 196150 97020 196350 97090
rect 196650 97020 196850 97090
rect 197150 97020 197350 97090
rect 197650 97020 197850 97090
rect 198150 97020 198350 97090
rect 198650 97020 198850 97090
rect 199150 97020 199350 97090
rect 199650 97020 199850 97090
rect 200150 97020 200350 97090
rect 200650 97020 200850 97090
rect 201150 97020 201350 97090
rect 201650 97020 201850 97090
rect 202150 97020 202350 97090
rect 202650 97020 202850 97090
rect 203150 97020 203350 97090
rect 203650 97020 203850 97090
rect 204150 97020 204350 97090
rect 204650 97020 204850 97090
rect 205150 97020 205350 97090
rect 205650 97020 205850 97090
rect 206150 97020 206350 97090
rect 206650 97020 206850 97090
rect 207150 97020 207350 97090
rect 207650 97020 207850 97090
rect 196150 96910 196350 96980
rect 196650 96910 196850 96980
rect 197150 96910 197350 96980
rect 197650 96910 197850 96980
rect 198150 96910 198350 96980
rect 198650 96910 198850 96980
rect 199150 96910 199350 96980
rect 199650 96910 199850 96980
rect 200150 96910 200350 96980
rect 200650 96910 200850 96980
rect 201150 96910 201350 96980
rect 201650 96910 201850 96980
rect 202150 96910 202350 96980
rect 202650 96910 202850 96980
rect 203150 96910 203350 96980
rect 203650 96910 203850 96980
rect 204150 96910 204350 96980
rect 204650 96910 204850 96980
rect 205150 96910 205350 96980
rect 205650 96910 205850 96980
rect 206150 96910 206350 96980
rect 206650 96910 206850 96980
rect 207150 96910 207350 96980
rect 207650 96910 207850 96980
rect 196020 96650 196090 96850
rect 196410 96650 196480 96850
rect 196520 96650 196590 96850
rect 196910 96650 196980 96850
rect 197020 96650 197090 96850
rect 197410 96650 197480 96850
rect 197520 96650 197590 96850
rect 197910 96650 197980 96850
rect 198020 96650 198090 96850
rect 198410 96650 198480 96850
rect 198520 96650 198590 96850
rect 198910 96650 198980 96850
rect 199020 96650 199090 96850
rect 199410 96650 199480 96850
rect 199520 96650 199590 96850
rect 199910 96650 199980 96850
rect 200020 96650 200090 96850
rect 200410 96650 200480 96850
rect 200520 96650 200590 96850
rect 200910 96650 200980 96850
rect 201020 96650 201090 96850
rect 201410 96650 201480 96850
rect 201520 96650 201590 96850
rect 201910 96650 201980 96850
rect 202020 96650 202090 96850
rect 202410 96650 202480 96850
rect 202520 96650 202590 96850
rect 202910 96650 202980 96850
rect 203020 96650 203090 96850
rect 203410 96650 203480 96850
rect 203520 96650 203590 96850
rect 203910 96650 203980 96850
rect 204020 96650 204090 96850
rect 204410 96650 204480 96850
rect 204520 96650 204590 96850
rect 204910 96650 204980 96850
rect 205020 96650 205090 96850
rect 205410 96650 205480 96850
rect 205520 96650 205590 96850
rect 205910 96650 205980 96850
rect 206020 96650 206090 96850
rect 206410 96650 206480 96850
rect 206520 96650 206590 96850
rect 206910 96650 206980 96850
rect 207020 96650 207090 96850
rect 207410 96650 207480 96850
rect 207520 96650 207590 96850
rect 207910 96650 207980 96850
rect 196150 96520 196350 96590
rect 196650 96520 196850 96590
rect 197150 96520 197350 96590
rect 197650 96520 197850 96590
rect 198150 96520 198350 96590
rect 198650 96520 198850 96590
rect 199150 96520 199350 96590
rect 199650 96520 199850 96590
rect 200150 96520 200350 96590
rect 200650 96520 200850 96590
rect 201150 96520 201350 96590
rect 201650 96520 201850 96590
rect 202150 96520 202350 96590
rect 202650 96520 202850 96590
rect 203150 96520 203350 96590
rect 203650 96520 203850 96590
rect 204150 96520 204350 96590
rect 204650 96520 204850 96590
rect 205150 96520 205350 96590
rect 205650 96520 205850 96590
rect 206150 96520 206350 96590
rect 206650 96520 206850 96590
rect 207150 96520 207350 96590
rect 207650 96520 207850 96590
rect 196150 96410 196350 96480
rect 196650 96410 196850 96480
rect 197150 96410 197350 96480
rect 197650 96410 197850 96480
rect 198150 96410 198350 96480
rect 198650 96410 198850 96480
rect 199150 96410 199350 96480
rect 199650 96410 199850 96480
rect 200150 96410 200350 96480
rect 200650 96410 200850 96480
rect 201150 96410 201350 96480
rect 201650 96410 201850 96480
rect 202150 96410 202350 96480
rect 202650 96410 202850 96480
rect 203150 96410 203350 96480
rect 203650 96410 203850 96480
rect 204150 96410 204350 96480
rect 204650 96410 204850 96480
rect 205150 96410 205350 96480
rect 205650 96410 205850 96480
rect 206150 96410 206350 96480
rect 206650 96410 206850 96480
rect 207150 96410 207350 96480
rect 207650 96410 207850 96480
rect 196020 96150 196090 96350
rect 196410 96150 196480 96350
rect 196520 96150 196590 96350
rect 196910 96150 196980 96350
rect 197020 96150 197090 96350
rect 197410 96150 197480 96350
rect 197520 96150 197590 96350
rect 197910 96150 197980 96350
rect 198020 96150 198090 96350
rect 198410 96150 198480 96350
rect 198520 96150 198590 96350
rect 198910 96150 198980 96350
rect 199020 96150 199090 96350
rect 199410 96150 199480 96350
rect 199520 96150 199590 96350
rect 199910 96150 199980 96350
rect 200020 96150 200090 96350
rect 200410 96150 200480 96350
rect 200520 96150 200590 96350
rect 200910 96150 200980 96350
rect 201020 96150 201090 96350
rect 201410 96150 201480 96350
rect 201520 96150 201590 96350
rect 201910 96150 201980 96350
rect 202020 96150 202090 96350
rect 202410 96150 202480 96350
rect 202520 96150 202590 96350
rect 202910 96150 202980 96350
rect 203020 96150 203090 96350
rect 203410 96150 203480 96350
rect 203520 96150 203590 96350
rect 203910 96150 203980 96350
rect 204020 96150 204090 96350
rect 204410 96150 204480 96350
rect 204520 96150 204590 96350
rect 204910 96150 204980 96350
rect 205020 96150 205090 96350
rect 205410 96150 205480 96350
rect 205520 96150 205590 96350
rect 205910 96150 205980 96350
rect 206020 96150 206090 96350
rect 206410 96150 206480 96350
rect 206520 96150 206590 96350
rect 206910 96150 206980 96350
rect 207020 96150 207090 96350
rect 207410 96150 207480 96350
rect 207520 96150 207590 96350
rect 207910 96150 207980 96350
rect 196150 96020 196350 96090
rect 196650 96020 196850 96090
rect 197150 96020 197350 96090
rect 197650 96020 197850 96090
rect 198150 96020 198350 96090
rect 198650 96020 198850 96090
rect 199150 96020 199350 96090
rect 199650 96020 199850 96090
rect 200150 96020 200350 96090
rect 200650 96020 200850 96090
rect 201150 96020 201350 96090
rect 201650 96020 201850 96090
rect 202150 96020 202350 96090
rect 202650 96020 202850 96090
rect 203150 96020 203350 96090
rect 203650 96020 203850 96090
rect 204150 96020 204350 96090
rect 204650 96020 204850 96090
rect 205150 96020 205350 96090
rect 205650 96020 205850 96090
rect 206150 96020 206350 96090
rect 206650 96020 206850 96090
rect 207150 96020 207350 96090
rect 207650 96020 207850 96090
rect 196150 95910 196350 95980
rect 196650 95910 196850 95980
rect 197150 95910 197350 95980
rect 197650 95910 197850 95980
rect 198150 95910 198350 95980
rect 198650 95910 198850 95980
rect 199150 95910 199350 95980
rect 199650 95910 199850 95980
rect 200150 95910 200350 95980
rect 200650 95910 200850 95980
rect 201150 95910 201350 95980
rect 201650 95910 201850 95980
rect 202150 95910 202350 95980
rect 202650 95910 202850 95980
rect 203150 95910 203350 95980
rect 203650 95910 203850 95980
rect 204150 95910 204350 95980
rect 204650 95910 204850 95980
rect 205150 95910 205350 95980
rect 205650 95910 205850 95980
rect 206150 95910 206350 95980
rect 206650 95910 206850 95980
rect 207150 95910 207350 95980
rect 207650 95910 207850 95980
rect 196020 95650 196090 95850
rect 196410 95650 196480 95850
rect 196520 95650 196590 95850
rect 196910 95650 196980 95850
rect 197020 95650 197090 95850
rect 197410 95650 197480 95850
rect 197520 95650 197590 95850
rect 197910 95650 197980 95850
rect 198020 95650 198090 95850
rect 198410 95650 198480 95850
rect 198520 95650 198590 95850
rect 198910 95650 198980 95850
rect 199020 95650 199090 95850
rect 199410 95650 199480 95850
rect 199520 95650 199590 95850
rect 199910 95650 199980 95850
rect 200020 95650 200090 95850
rect 200410 95650 200480 95850
rect 200520 95650 200590 95850
rect 200910 95650 200980 95850
rect 201020 95650 201090 95850
rect 201410 95650 201480 95850
rect 201520 95650 201590 95850
rect 201910 95650 201980 95850
rect 202020 95650 202090 95850
rect 202410 95650 202480 95850
rect 202520 95650 202590 95850
rect 202910 95650 202980 95850
rect 203020 95650 203090 95850
rect 203410 95650 203480 95850
rect 203520 95650 203590 95850
rect 203910 95650 203980 95850
rect 204020 95650 204090 95850
rect 204410 95650 204480 95850
rect 204520 95650 204590 95850
rect 204910 95650 204980 95850
rect 205020 95650 205090 95850
rect 205410 95650 205480 95850
rect 205520 95650 205590 95850
rect 205910 95650 205980 95850
rect 206020 95650 206090 95850
rect 206410 95650 206480 95850
rect 206520 95650 206590 95850
rect 206910 95650 206980 95850
rect 207020 95650 207090 95850
rect 207410 95650 207480 95850
rect 207520 95650 207590 95850
rect 207910 95650 207980 95850
rect 196150 95520 196350 95590
rect 196650 95520 196850 95590
rect 197150 95520 197350 95590
rect 197650 95520 197850 95590
rect 198150 95520 198350 95590
rect 198650 95520 198850 95590
rect 199150 95520 199350 95590
rect 199650 95520 199850 95590
rect 200150 95520 200350 95590
rect 200650 95520 200850 95590
rect 201150 95520 201350 95590
rect 201650 95520 201850 95590
rect 202150 95520 202350 95590
rect 202650 95520 202850 95590
rect 203150 95520 203350 95590
rect 203650 95520 203850 95590
rect 204150 95520 204350 95590
rect 204650 95520 204850 95590
rect 205150 95520 205350 95590
rect 205650 95520 205850 95590
rect 206150 95520 206350 95590
rect 206650 95520 206850 95590
rect 207150 95520 207350 95590
rect 207650 95520 207850 95590
rect 196150 95410 196350 95480
rect 196650 95410 196850 95480
rect 197150 95410 197350 95480
rect 197650 95410 197850 95480
rect 198150 95410 198350 95480
rect 198650 95410 198850 95480
rect 199150 95410 199350 95480
rect 199650 95410 199850 95480
rect 200150 95410 200350 95480
rect 200650 95410 200850 95480
rect 201150 95410 201350 95480
rect 201650 95410 201850 95480
rect 202150 95410 202350 95480
rect 202650 95410 202850 95480
rect 203150 95410 203350 95480
rect 203650 95410 203850 95480
rect 204150 95410 204350 95480
rect 204650 95410 204850 95480
rect 205150 95410 205350 95480
rect 205650 95410 205850 95480
rect 206150 95410 206350 95480
rect 206650 95410 206850 95480
rect 207150 95410 207350 95480
rect 207650 95410 207850 95480
rect 196020 95150 196090 95350
rect 196410 95150 196480 95350
rect 196520 95150 196590 95350
rect 196910 95150 196980 95350
rect 197020 95150 197090 95350
rect 197410 95150 197480 95350
rect 197520 95150 197590 95350
rect 197910 95150 197980 95350
rect 198020 95150 198090 95350
rect 198410 95150 198480 95350
rect 198520 95150 198590 95350
rect 198910 95150 198980 95350
rect 199020 95150 199090 95350
rect 199410 95150 199480 95350
rect 199520 95150 199590 95350
rect 199910 95150 199980 95350
rect 200020 95150 200090 95350
rect 200410 95150 200480 95350
rect 200520 95150 200590 95350
rect 200910 95150 200980 95350
rect 201020 95150 201090 95350
rect 201410 95150 201480 95350
rect 201520 95150 201590 95350
rect 201910 95150 201980 95350
rect 202020 95150 202090 95350
rect 202410 95150 202480 95350
rect 202520 95150 202590 95350
rect 202910 95150 202980 95350
rect 203020 95150 203090 95350
rect 203410 95150 203480 95350
rect 203520 95150 203590 95350
rect 203910 95150 203980 95350
rect 204020 95150 204090 95350
rect 204410 95150 204480 95350
rect 204520 95150 204590 95350
rect 204910 95150 204980 95350
rect 205020 95150 205090 95350
rect 205410 95150 205480 95350
rect 205520 95150 205590 95350
rect 205910 95150 205980 95350
rect 206020 95150 206090 95350
rect 206410 95150 206480 95350
rect 206520 95150 206590 95350
rect 206910 95150 206980 95350
rect 207020 95150 207090 95350
rect 207410 95150 207480 95350
rect 207520 95150 207590 95350
rect 207910 95150 207980 95350
rect 196150 95020 196350 95090
rect 196650 95020 196850 95090
rect 197150 95020 197350 95090
rect 197650 95020 197850 95090
rect 198150 95020 198350 95090
rect 198650 95020 198850 95090
rect 199150 95020 199350 95090
rect 199650 95020 199850 95090
rect 200150 95020 200350 95090
rect 200650 95020 200850 95090
rect 201150 95020 201350 95090
rect 201650 95020 201850 95090
rect 202150 95020 202350 95090
rect 202650 95020 202850 95090
rect 203150 95020 203350 95090
rect 203650 95020 203850 95090
rect 204150 95020 204350 95090
rect 204650 95020 204850 95090
rect 205150 95020 205350 95090
rect 205650 95020 205850 95090
rect 206150 95020 206350 95090
rect 206650 95020 206850 95090
rect 207150 95020 207350 95090
rect 207650 95020 207850 95090
rect 196150 94910 196350 94980
rect 196650 94910 196850 94980
rect 197150 94910 197350 94980
rect 197650 94910 197850 94980
rect 198150 94910 198350 94980
rect 198650 94910 198850 94980
rect 199150 94910 199350 94980
rect 199650 94910 199850 94980
rect 200150 94910 200350 94980
rect 200650 94910 200850 94980
rect 201150 94910 201350 94980
rect 201650 94910 201850 94980
rect 202150 94910 202350 94980
rect 202650 94910 202850 94980
rect 203150 94910 203350 94980
rect 203650 94910 203850 94980
rect 204150 94910 204350 94980
rect 204650 94910 204850 94980
rect 205150 94910 205350 94980
rect 205650 94910 205850 94980
rect 206150 94910 206350 94980
rect 206650 94910 206850 94980
rect 207150 94910 207350 94980
rect 207650 94910 207850 94980
rect 196020 94650 196090 94850
rect 196410 94650 196480 94850
rect 196520 94650 196590 94850
rect 196910 94650 196980 94850
rect 197020 94650 197090 94850
rect 197410 94650 197480 94850
rect 197520 94650 197590 94850
rect 197910 94650 197980 94850
rect 198020 94650 198090 94850
rect 198410 94650 198480 94850
rect 198520 94650 198590 94850
rect 198910 94650 198980 94850
rect 199020 94650 199090 94850
rect 199410 94650 199480 94850
rect 199520 94650 199590 94850
rect 199910 94650 199980 94850
rect 200020 94650 200090 94850
rect 200410 94650 200480 94850
rect 200520 94650 200590 94850
rect 200910 94650 200980 94850
rect 201020 94650 201090 94850
rect 201410 94650 201480 94850
rect 201520 94650 201590 94850
rect 201910 94650 201980 94850
rect 202020 94650 202090 94850
rect 202410 94650 202480 94850
rect 202520 94650 202590 94850
rect 202910 94650 202980 94850
rect 203020 94650 203090 94850
rect 203410 94650 203480 94850
rect 203520 94650 203590 94850
rect 203910 94650 203980 94850
rect 204020 94650 204090 94850
rect 204410 94650 204480 94850
rect 204520 94650 204590 94850
rect 204910 94650 204980 94850
rect 205020 94650 205090 94850
rect 205410 94650 205480 94850
rect 205520 94650 205590 94850
rect 205910 94650 205980 94850
rect 206020 94650 206090 94850
rect 206410 94650 206480 94850
rect 206520 94650 206590 94850
rect 206910 94650 206980 94850
rect 207020 94650 207090 94850
rect 207410 94650 207480 94850
rect 207520 94650 207590 94850
rect 207910 94650 207980 94850
rect 196150 94520 196350 94590
rect 196650 94520 196850 94590
rect 197150 94520 197350 94590
rect 197650 94520 197850 94590
rect 198150 94520 198350 94590
rect 198650 94520 198850 94590
rect 199150 94520 199350 94590
rect 199650 94520 199850 94590
rect 200150 94520 200350 94590
rect 200650 94520 200850 94590
rect 201150 94520 201350 94590
rect 201650 94520 201850 94590
rect 202150 94520 202350 94590
rect 202650 94520 202850 94590
rect 203150 94520 203350 94590
rect 203650 94520 203850 94590
rect 204150 94520 204350 94590
rect 204650 94520 204850 94590
rect 205150 94520 205350 94590
rect 205650 94520 205850 94590
rect 206150 94520 206350 94590
rect 206650 94520 206850 94590
rect 207150 94520 207350 94590
rect 207650 94520 207850 94590
rect 196150 94410 196350 94480
rect 196650 94410 196850 94480
rect 197150 94410 197350 94480
rect 197650 94410 197850 94480
rect 198150 94410 198350 94480
rect 198650 94410 198850 94480
rect 199150 94410 199350 94480
rect 199650 94410 199850 94480
rect 200150 94410 200350 94480
rect 200650 94410 200850 94480
rect 201150 94410 201350 94480
rect 201650 94410 201850 94480
rect 202150 94410 202350 94480
rect 202650 94410 202850 94480
rect 203150 94410 203350 94480
rect 203650 94410 203850 94480
rect 204150 94410 204350 94480
rect 204650 94410 204850 94480
rect 205150 94410 205350 94480
rect 205650 94410 205850 94480
rect 206150 94410 206350 94480
rect 206650 94410 206850 94480
rect 207150 94410 207350 94480
rect 207650 94410 207850 94480
rect 196020 94150 196090 94350
rect 196410 94150 196480 94350
rect 196520 94150 196590 94350
rect 196910 94150 196980 94350
rect 197020 94150 197090 94350
rect 197410 94150 197480 94350
rect 197520 94150 197590 94350
rect 197910 94150 197980 94350
rect 198020 94150 198090 94350
rect 198410 94150 198480 94350
rect 198520 94150 198590 94350
rect 198910 94150 198980 94350
rect 199020 94150 199090 94350
rect 199410 94150 199480 94350
rect 199520 94150 199590 94350
rect 199910 94150 199980 94350
rect 200020 94150 200090 94350
rect 200410 94150 200480 94350
rect 200520 94150 200590 94350
rect 200910 94150 200980 94350
rect 201020 94150 201090 94350
rect 201410 94150 201480 94350
rect 201520 94150 201590 94350
rect 201910 94150 201980 94350
rect 202020 94150 202090 94350
rect 202410 94150 202480 94350
rect 202520 94150 202590 94350
rect 202910 94150 202980 94350
rect 203020 94150 203090 94350
rect 203410 94150 203480 94350
rect 203520 94150 203590 94350
rect 203910 94150 203980 94350
rect 204020 94150 204090 94350
rect 204410 94150 204480 94350
rect 204520 94150 204590 94350
rect 204910 94150 204980 94350
rect 205020 94150 205090 94350
rect 205410 94150 205480 94350
rect 205520 94150 205590 94350
rect 205910 94150 205980 94350
rect 206020 94150 206090 94350
rect 206410 94150 206480 94350
rect 206520 94150 206590 94350
rect 206910 94150 206980 94350
rect 207020 94150 207090 94350
rect 207410 94150 207480 94350
rect 207520 94150 207590 94350
rect 207910 94150 207980 94350
rect 196150 94020 196350 94090
rect 196650 94020 196850 94090
rect 197150 94020 197350 94090
rect 197650 94020 197850 94090
rect 198150 94020 198350 94090
rect 198650 94020 198850 94090
rect 199150 94020 199350 94090
rect 199650 94020 199850 94090
rect 200150 94020 200350 94090
rect 200650 94020 200850 94090
rect 201150 94020 201350 94090
rect 201650 94020 201850 94090
rect 202150 94020 202350 94090
rect 202650 94020 202850 94090
rect 203150 94020 203350 94090
rect 203650 94020 203850 94090
rect 204150 94020 204350 94090
rect 204650 94020 204850 94090
rect 205150 94020 205350 94090
rect 205650 94020 205850 94090
rect 206150 94020 206350 94090
rect 206650 94020 206850 94090
rect 207150 94020 207350 94090
rect 207650 94020 207850 94090
rect 196150 93910 196350 93980
rect 196650 93910 196850 93980
rect 197150 93910 197350 93980
rect 197650 93910 197850 93980
rect 198150 93910 198350 93980
rect 198650 93910 198850 93980
rect 199150 93910 199350 93980
rect 199650 93910 199850 93980
rect 200150 93910 200350 93980
rect 200650 93910 200850 93980
rect 201150 93910 201350 93980
rect 201650 93910 201850 93980
rect 202150 93910 202350 93980
rect 202650 93910 202850 93980
rect 203150 93910 203350 93980
rect 203650 93910 203850 93980
rect 204150 93910 204350 93980
rect 204650 93910 204850 93980
rect 205150 93910 205350 93980
rect 205650 93910 205850 93980
rect 206150 93910 206350 93980
rect 206650 93910 206850 93980
rect 207150 93910 207350 93980
rect 207650 93910 207850 93980
rect 196020 93650 196090 93850
rect 196410 93650 196480 93850
rect 196520 93650 196590 93850
rect 196910 93650 196980 93850
rect 197020 93650 197090 93850
rect 197410 93650 197480 93850
rect 197520 93650 197590 93850
rect 197910 93650 197980 93850
rect 198020 93650 198090 93850
rect 198410 93650 198480 93850
rect 198520 93650 198590 93850
rect 198910 93650 198980 93850
rect 199020 93650 199090 93850
rect 199410 93650 199480 93850
rect 199520 93650 199590 93850
rect 199910 93650 199980 93850
rect 200020 93650 200090 93850
rect 200410 93650 200480 93850
rect 200520 93650 200590 93850
rect 200910 93650 200980 93850
rect 201020 93650 201090 93850
rect 201410 93650 201480 93850
rect 201520 93650 201590 93850
rect 201910 93650 201980 93850
rect 202020 93650 202090 93850
rect 202410 93650 202480 93850
rect 202520 93650 202590 93850
rect 202910 93650 202980 93850
rect 203020 93650 203090 93850
rect 203410 93650 203480 93850
rect 203520 93650 203590 93850
rect 203910 93650 203980 93850
rect 204020 93650 204090 93850
rect 204410 93650 204480 93850
rect 204520 93650 204590 93850
rect 204910 93650 204980 93850
rect 205020 93650 205090 93850
rect 205410 93650 205480 93850
rect 205520 93650 205590 93850
rect 205910 93650 205980 93850
rect 206020 93650 206090 93850
rect 206410 93650 206480 93850
rect 206520 93650 206590 93850
rect 206910 93650 206980 93850
rect 207020 93650 207090 93850
rect 207410 93650 207480 93850
rect 207520 93650 207590 93850
rect 207910 93650 207980 93850
rect 196150 93520 196350 93590
rect 196650 93520 196850 93590
rect 197150 93520 197350 93590
rect 197650 93520 197850 93590
rect 198150 93520 198350 93590
rect 198650 93520 198850 93590
rect 199150 93520 199350 93590
rect 199650 93520 199850 93590
rect 200150 93520 200350 93590
rect 200650 93520 200850 93590
rect 201150 93520 201350 93590
rect 201650 93520 201850 93590
rect 202150 93520 202350 93590
rect 202650 93520 202850 93590
rect 203150 93520 203350 93590
rect 203650 93520 203850 93590
rect 204150 93520 204350 93590
rect 204650 93520 204850 93590
rect 205150 93520 205350 93590
rect 205650 93520 205850 93590
rect 206150 93520 206350 93590
rect 206650 93520 206850 93590
rect 207150 93520 207350 93590
rect 207650 93520 207850 93590
rect 196150 93410 196350 93480
rect 196650 93410 196850 93480
rect 197150 93410 197350 93480
rect 197650 93410 197850 93480
rect 198150 93410 198350 93480
rect 198650 93410 198850 93480
rect 199150 93410 199350 93480
rect 199650 93410 199850 93480
rect 200150 93410 200350 93480
rect 200650 93410 200850 93480
rect 201150 93410 201350 93480
rect 201650 93410 201850 93480
rect 202150 93410 202350 93480
rect 202650 93410 202850 93480
rect 203150 93410 203350 93480
rect 203650 93410 203850 93480
rect 204150 93410 204350 93480
rect 204650 93410 204850 93480
rect 205150 93410 205350 93480
rect 205650 93410 205850 93480
rect 206150 93410 206350 93480
rect 206650 93410 206850 93480
rect 207150 93410 207350 93480
rect 207650 93410 207850 93480
rect 196020 93150 196090 93350
rect 196410 93150 196480 93350
rect 196520 93150 196590 93350
rect 196910 93150 196980 93350
rect 197020 93150 197090 93350
rect 197410 93150 197480 93350
rect 197520 93150 197590 93350
rect 197910 93150 197980 93350
rect 198020 93150 198090 93350
rect 198410 93150 198480 93350
rect 198520 93150 198590 93350
rect 198910 93150 198980 93350
rect 199020 93150 199090 93350
rect 199410 93150 199480 93350
rect 199520 93150 199590 93350
rect 199910 93150 199980 93350
rect 200020 93150 200090 93350
rect 200410 93150 200480 93350
rect 200520 93150 200590 93350
rect 200910 93150 200980 93350
rect 201020 93150 201090 93350
rect 201410 93150 201480 93350
rect 201520 93150 201590 93350
rect 201910 93150 201980 93350
rect 202020 93150 202090 93350
rect 202410 93150 202480 93350
rect 202520 93150 202590 93350
rect 202910 93150 202980 93350
rect 203020 93150 203090 93350
rect 203410 93150 203480 93350
rect 203520 93150 203590 93350
rect 203910 93150 203980 93350
rect 204020 93150 204090 93350
rect 204410 93150 204480 93350
rect 204520 93150 204590 93350
rect 204910 93150 204980 93350
rect 205020 93150 205090 93350
rect 205410 93150 205480 93350
rect 205520 93150 205590 93350
rect 205910 93150 205980 93350
rect 206020 93150 206090 93350
rect 206410 93150 206480 93350
rect 206520 93150 206590 93350
rect 206910 93150 206980 93350
rect 207020 93150 207090 93350
rect 207410 93150 207480 93350
rect 207520 93150 207590 93350
rect 207910 93150 207980 93350
rect 196150 93020 196350 93090
rect 196650 93020 196850 93090
rect 197150 93020 197350 93090
rect 197650 93020 197850 93090
rect 198150 93020 198350 93090
rect 198650 93020 198850 93090
rect 199150 93020 199350 93090
rect 199650 93020 199850 93090
rect 200150 93020 200350 93090
rect 200650 93020 200850 93090
rect 201150 93020 201350 93090
rect 201650 93020 201850 93090
rect 202150 93020 202350 93090
rect 202650 93020 202850 93090
rect 203150 93020 203350 93090
rect 203650 93020 203850 93090
rect 204150 93020 204350 93090
rect 204650 93020 204850 93090
rect 205150 93020 205350 93090
rect 205650 93020 205850 93090
rect 206150 93020 206350 93090
rect 206650 93020 206850 93090
rect 207150 93020 207350 93090
rect 207650 93020 207850 93090
rect 196150 92910 196350 92980
rect 196650 92910 196850 92980
rect 197150 92910 197350 92980
rect 197650 92910 197850 92980
rect 198150 92910 198350 92980
rect 198650 92910 198850 92980
rect 199150 92910 199350 92980
rect 199650 92910 199850 92980
rect 200150 92910 200350 92980
rect 200650 92910 200850 92980
rect 201150 92910 201350 92980
rect 201650 92910 201850 92980
rect 202150 92910 202350 92980
rect 202650 92910 202850 92980
rect 203150 92910 203350 92980
rect 203650 92910 203850 92980
rect 204150 92910 204350 92980
rect 204650 92910 204850 92980
rect 205150 92910 205350 92980
rect 205650 92910 205850 92980
rect 206150 92910 206350 92980
rect 206650 92910 206850 92980
rect 207150 92910 207350 92980
rect 207650 92910 207850 92980
rect 196020 92650 196090 92850
rect 196410 92650 196480 92850
rect 196520 92650 196590 92850
rect 196910 92650 196980 92850
rect 197020 92650 197090 92850
rect 197410 92650 197480 92850
rect 197520 92650 197590 92850
rect 197910 92650 197980 92850
rect 198020 92650 198090 92850
rect 198410 92650 198480 92850
rect 198520 92650 198590 92850
rect 198910 92650 198980 92850
rect 199020 92650 199090 92850
rect 199410 92650 199480 92850
rect 199520 92650 199590 92850
rect 199910 92650 199980 92850
rect 200020 92650 200090 92850
rect 200410 92650 200480 92850
rect 200520 92650 200590 92850
rect 200910 92650 200980 92850
rect 201020 92650 201090 92850
rect 201410 92650 201480 92850
rect 201520 92650 201590 92850
rect 201910 92650 201980 92850
rect 202020 92650 202090 92850
rect 202410 92650 202480 92850
rect 202520 92650 202590 92850
rect 202910 92650 202980 92850
rect 203020 92650 203090 92850
rect 203410 92650 203480 92850
rect 203520 92650 203590 92850
rect 203910 92650 203980 92850
rect 204020 92650 204090 92850
rect 204410 92650 204480 92850
rect 204520 92650 204590 92850
rect 204910 92650 204980 92850
rect 205020 92650 205090 92850
rect 205410 92650 205480 92850
rect 205520 92650 205590 92850
rect 205910 92650 205980 92850
rect 206020 92650 206090 92850
rect 206410 92650 206480 92850
rect 206520 92650 206590 92850
rect 206910 92650 206980 92850
rect 207020 92650 207090 92850
rect 207410 92650 207480 92850
rect 207520 92650 207590 92850
rect 207910 92650 207980 92850
rect 196150 92520 196350 92590
rect 196650 92520 196850 92590
rect 197150 92520 197350 92590
rect 197650 92520 197850 92590
rect 198150 92520 198350 92590
rect 198650 92520 198850 92590
rect 199150 92520 199350 92590
rect 199650 92520 199850 92590
rect 200150 92520 200350 92590
rect 200650 92520 200850 92590
rect 201150 92520 201350 92590
rect 201650 92520 201850 92590
rect 202150 92520 202350 92590
rect 202650 92520 202850 92590
rect 203150 92520 203350 92590
rect 203650 92520 203850 92590
rect 204150 92520 204350 92590
rect 204650 92520 204850 92590
rect 205150 92520 205350 92590
rect 205650 92520 205850 92590
rect 206150 92520 206350 92590
rect 206650 92520 206850 92590
rect 207150 92520 207350 92590
rect 207650 92520 207850 92590
rect 196150 92410 196350 92480
rect 196650 92410 196850 92480
rect 197150 92410 197350 92480
rect 197650 92410 197850 92480
rect 198150 92410 198350 92480
rect 198650 92410 198850 92480
rect 199150 92410 199350 92480
rect 199650 92410 199850 92480
rect 200150 92410 200350 92480
rect 200650 92410 200850 92480
rect 201150 92410 201350 92480
rect 201650 92410 201850 92480
rect 202150 92410 202350 92480
rect 202650 92410 202850 92480
rect 203150 92410 203350 92480
rect 203650 92410 203850 92480
rect 204150 92410 204350 92480
rect 204650 92410 204850 92480
rect 205150 92410 205350 92480
rect 205650 92410 205850 92480
rect 206150 92410 206350 92480
rect 206650 92410 206850 92480
rect 207150 92410 207350 92480
rect 207650 92410 207850 92480
rect 196020 92150 196090 92350
rect 196410 92150 196480 92350
rect 196520 92150 196590 92350
rect 196910 92150 196980 92350
rect 197020 92150 197090 92350
rect 197410 92150 197480 92350
rect 197520 92150 197590 92350
rect 197910 92150 197980 92350
rect 198020 92150 198090 92350
rect 198410 92150 198480 92350
rect 198520 92150 198590 92350
rect 198910 92150 198980 92350
rect 199020 92150 199090 92350
rect 199410 92150 199480 92350
rect 199520 92150 199590 92350
rect 199910 92150 199980 92350
rect 200020 92150 200090 92350
rect 200410 92150 200480 92350
rect 200520 92150 200590 92350
rect 200910 92150 200980 92350
rect 201020 92150 201090 92350
rect 201410 92150 201480 92350
rect 201520 92150 201590 92350
rect 201910 92150 201980 92350
rect 202020 92150 202090 92350
rect 202410 92150 202480 92350
rect 202520 92150 202590 92350
rect 202910 92150 202980 92350
rect 203020 92150 203090 92350
rect 203410 92150 203480 92350
rect 203520 92150 203590 92350
rect 203910 92150 203980 92350
rect 204020 92150 204090 92350
rect 204410 92150 204480 92350
rect 204520 92150 204590 92350
rect 204910 92150 204980 92350
rect 205020 92150 205090 92350
rect 205410 92150 205480 92350
rect 205520 92150 205590 92350
rect 205910 92150 205980 92350
rect 206020 92150 206090 92350
rect 206410 92150 206480 92350
rect 206520 92150 206590 92350
rect 206910 92150 206980 92350
rect 207020 92150 207090 92350
rect 207410 92150 207480 92350
rect 207520 92150 207590 92350
rect 207910 92150 207980 92350
rect 196150 92020 196350 92090
rect 196650 92020 196850 92090
rect 197150 92020 197350 92090
rect 197650 92020 197850 92090
rect 198150 92020 198350 92090
rect 198650 92020 198850 92090
rect 199150 92020 199350 92090
rect 199650 92020 199850 92090
rect 200150 92020 200350 92090
rect 200650 92020 200850 92090
rect 201150 92020 201350 92090
rect 201650 92020 201850 92090
rect 202150 92020 202350 92090
rect 202650 92020 202850 92090
rect 203150 92020 203350 92090
rect 203650 92020 203850 92090
rect 204150 92020 204350 92090
rect 204650 92020 204850 92090
rect 205150 92020 205350 92090
rect 205650 92020 205850 92090
rect 206150 92020 206350 92090
rect 206650 92020 206850 92090
rect 207150 92020 207350 92090
rect 207650 92020 207850 92090
rect 196150 91910 196350 91980
rect 196650 91910 196850 91980
rect 197150 91910 197350 91980
rect 197650 91910 197850 91980
rect 198150 91910 198350 91980
rect 198650 91910 198850 91980
rect 199150 91910 199350 91980
rect 199650 91910 199850 91980
rect 200150 91910 200350 91980
rect 200650 91910 200850 91980
rect 201150 91910 201350 91980
rect 201650 91910 201850 91980
rect 202150 91910 202350 91980
rect 202650 91910 202850 91980
rect 203150 91910 203350 91980
rect 203650 91910 203850 91980
rect 204150 91910 204350 91980
rect 204650 91910 204850 91980
rect 205150 91910 205350 91980
rect 205650 91910 205850 91980
rect 206150 91910 206350 91980
rect 206650 91910 206850 91980
rect 207150 91910 207350 91980
rect 207650 91910 207850 91980
rect 196020 91650 196090 91850
rect 196410 91650 196480 91850
rect 196520 91650 196590 91850
rect 196910 91650 196980 91850
rect 197020 91650 197090 91850
rect 197410 91650 197480 91850
rect 197520 91650 197590 91850
rect 197910 91650 197980 91850
rect 198020 91650 198090 91850
rect 198410 91650 198480 91850
rect 198520 91650 198590 91850
rect 198910 91650 198980 91850
rect 199020 91650 199090 91850
rect 199410 91650 199480 91850
rect 199520 91650 199590 91850
rect 199910 91650 199980 91850
rect 200020 91650 200090 91850
rect 200410 91650 200480 91850
rect 200520 91650 200590 91850
rect 200910 91650 200980 91850
rect 201020 91650 201090 91850
rect 201410 91650 201480 91850
rect 201520 91650 201590 91850
rect 201910 91650 201980 91850
rect 202020 91650 202090 91850
rect 202410 91650 202480 91850
rect 202520 91650 202590 91850
rect 202910 91650 202980 91850
rect 203020 91650 203090 91850
rect 203410 91650 203480 91850
rect 203520 91650 203590 91850
rect 203910 91650 203980 91850
rect 204020 91650 204090 91850
rect 204410 91650 204480 91850
rect 204520 91650 204590 91850
rect 204910 91650 204980 91850
rect 205020 91650 205090 91850
rect 205410 91650 205480 91850
rect 205520 91650 205590 91850
rect 205910 91650 205980 91850
rect 206020 91650 206090 91850
rect 206410 91650 206480 91850
rect 206520 91650 206590 91850
rect 206910 91650 206980 91850
rect 207020 91650 207090 91850
rect 207410 91650 207480 91850
rect 207520 91650 207590 91850
rect 207910 91650 207980 91850
rect 196150 91520 196350 91590
rect 196650 91520 196850 91590
rect 197150 91520 197350 91590
rect 197650 91520 197850 91590
rect 198150 91520 198350 91590
rect 198650 91520 198850 91590
rect 199150 91520 199350 91590
rect 199650 91520 199850 91590
rect 200150 91520 200350 91590
rect 200650 91520 200850 91590
rect 201150 91520 201350 91590
rect 201650 91520 201850 91590
rect 202150 91520 202350 91590
rect 202650 91520 202850 91590
rect 203150 91520 203350 91590
rect 203650 91520 203850 91590
rect 204150 91520 204350 91590
rect 204650 91520 204850 91590
rect 205150 91520 205350 91590
rect 205650 91520 205850 91590
rect 206150 91520 206350 91590
rect 206650 91520 206850 91590
rect 207150 91520 207350 91590
rect 207650 91520 207850 91590
rect 196150 91410 196350 91480
rect 196650 91410 196850 91480
rect 197150 91410 197350 91480
rect 197650 91410 197850 91480
rect 198150 91410 198350 91480
rect 198650 91410 198850 91480
rect 199150 91410 199350 91480
rect 199650 91410 199850 91480
rect 200150 91410 200350 91480
rect 200650 91410 200850 91480
rect 201150 91410 201350 91480
rect 201650 91410 201850 91480
rect 202150 91410 202350 91480
rect 202650 91410 202850 91480
rect 203150 91410 203350 91480
rect 203650 91410 203850 91480
rect 204150 91410 204350 91480
rect 204650 91410 204850 91480
rect 205150 91410 205350 91480
rect 205650 91410 205850 91480
rect 206150 91410 206350 91480
rect 206650 91410 206850 91480
rect 207150 91410 207350 91480
rect 207650 91410 207850 91480
rect 196020 91150 196090 91350
rect 196410 91150 196480 91350
rect 196520 91150 196590 91350
rect 196910 91150 196980 91350
rect 197020 91150 197090 91350
rect 197410 91150 197480 91350
rect 197520 91150 197590 91350
rect 197910 91150 197980 91350
rect 198020 91150 198090 91350
rect 198410 91150 198480 91350
rect 198520 91150 198590 91350
rect 198910 91150 198980 91350
rect 199020 91150 199090 91350
rect 199410 91150 199480 91350
rect 199520 91150 199590 91350
rect 199910 91150 199980 91350
rect 200020 91150 200090 91350
rect 200410 91150 200480 91350
rect 200520 91150 200590 91350
rect 200910 91150 200980 91350
rect 201020 91150 201090 91350
rect 201410 91150 201480 91350
rect 201520 91150 201590 91350
rect 201910 91150 201980 91350
rect 202020 91150 202090 91350
rect 202410 91150 202480 91350
rect 202520 91150 202590 91350
rect 202910 91150 202980 91350
rect 203020 91150 203090 91350
rect 203410 91150 203480 91350
rect 203520 91150 203590 91350
rect 203910 91150 203980 91350
rect 204020 91150 204090 91350
rect 204410 91150 204480 91350
rect 204520 91150 204590 91350
rect 204910 91150 204980 91350
rect 205020 91150 205090 91350
rect 205410 91150 205480 91350
rect 205520 91150 205590 91350
rect 205910 91150 205980 91350
rect 206020 91150 206090 91350
rect 206410 91150 206480 91350
rect 206520 91150 206590 91350
rect 206910 91150 206980 91350
rect 207020 91150 207090 91350
rect 207410 91150 207480 91350
rect 207520 91150 207590 91350
rect 207910 91150 207980 91350
rect 196150 91020 196350 91090
rect 196650 91020 196850 91090
rect 197150 91020 197350 91090
rect 197650 91020 197850 91090
rect 198150 91020 198350 91090
rect 198650 91020 198850 91090
rect 199150 91020 199350 91090
rect 199650 91020 199850 91090
rect 200150 91020 200350 91090
rect 200650 91020 200850 91090
rect 201150 91020 201350 91090
rect 201650 91020 201850 91090
rect 202150 91020 202350 91090
rect 202650 91020 202850 91090
rect 203150 91020 203350 91090
rect 203650 91020 203850 91090
rect 204150 91020 204350 91090
rect 204650 91020 204850 91090
rect 205150 91020 205350 91090
rect 205650 91020 205850 91090
rect 206150 91020 206350 91090
rect 206650 91020 206850 91090
rect 207150 91020 207350 91090
rect 207650 91020 207850 91090
rect 196150 90910 196350 90980
rect 196650 90910 196850 90980
rect 197150 90910 197350 90980
rect 197650 90910 197850 90980
rect 198150 90910 198350 90980
rect 198650 90910 198850 90980
rect 199150 90910 199350 90980
rect 199650 90910 199850 90980
rect 200150 90910 200350 90980
rect 200650 90910 200850 90980
rect 201150 90910 201350 90980
rect 201650 90910 201850 90980
rect 202150 90910 202350 90980
rect 202650 90910 202850 90980
rect 203150 90910 203350 90980
rect 203650 90910 203850 90980
rect 204150 90910 204350 90980
rect 204650 90910 204850 90980
rect 205150 90910 205350 90980
rect 205650 90910 205850 90980
rect 206150 90910 206350 90980
rect 206650 90910 206850 90980
rect 207150 90910 207350 90980
rect 207650 90910 207850 90980
rect 196020 90650 196090 90850
rect 196410 90650 196480 90850
rect 196520 90650 196590 90850
rect 196910 90650 196980 90850
rect 197020 90650 197090 90850
rect 197410 90650 197480 90850
rect 197520 90650 197590 90850
rect 197910 90650 197980 90850
rect 198020 90650 198090 90850
rect 198410 90650 198480 90850
rect 198520 90650 198590 90850
rect 198910 90650 198980 90850
rect 199020 90650 199090 90850
rect 199410 90650 199480 90850
rect 199520 90650 199590 90850
rect 199910 90650 199980 90850
rect 200020 90650 200090 90850
rect 200410 90650 200480 90850
rect 200520 90650 200590 90850
rect 200910 90650 200980 90850
rect 201020 90650 201090 90850
rect 201410 90650 201480 90850
rect 201520 90650 201590 90850
rect 201910 90650 201980 90850
rect 202020 90650 202090 90850
rect 202410 90650 202480 90850
rect 202520 90650 202590 90850
rect 202910 90650 202980 90850
rect 203020 90650 203090 90850
rect 203410 90650 203480 90850
rect 203520 90650 203590 90850
rect 203910 90650 203980 90850
rect 204020 90650 204090 90850
rect 204410 90650 204480 90850
rect 204520 90650 204590 90850
rect 204910 90650 204980 90850
rect 205020 90650 205090 90850
rect 205410 90650 205480 90850
rect 205520 90650 205590 90850
rect 205910 90650 205980 90850
rect 206020 90650 206090 90850
rect 206410 90650 206480 90850
rect 206520 90650 206590 90850
rect 206910 90650 206980 90850
rect 207020 90650 207090 90850
rect 207410 90650 207480 90850
rect 207520 90650 207590 90850
rect 207910 90650 207980 90850
rect 196150 90520 196350 90590
rect 196650 90520 196850 90590
rect 197150 90520 197350 90590
rect 197650 90520 197850 90590
rect 198150 90520 198350 90590
rect 198650 90520 198850 90590
rect 199150 90520 199350 90590
rect 199650 90520 199850 90590
rect 200150 90520 200350 90590
rect 200650 90520 200850 90590
rect 201150 90520 201350 90590
rect 201650 90520 201850 90590
rect 202150 90520 202350 90590
rect 202650 90520 202850 90590
rect 203150 90520 203350 90590
rect 203650 90520 203850 90590
rect 204150 90520 204350 90590
rect 204650 90520 204850 90590
rect 205150 90520 205350 90590
rect 205650 90520 205850 90590
rect 206150 90520 206350 90590
rect 206650 90520 206850 90590
rect 207150 90520 207350 90590
rect 207650 90520 207850 90590
rect 196150 90410 196350 90480
rect 196650 90410 196850 90480
rect 197150 90410 197350 90480
rect 197650 90410 197850 90480
rect 198150 90410 198350 90480
rect 198650 90410 198850 90480
rect 199150 90410 199350 90480
rect 199650 90410 199850 90480
rect 200150 90410 200350 90480
rect 200650 90410 200850 90480
rect 201150 90410 201350 90480
rect 201650 90410 201850 90480
rect 202150 90410 202350 90480
rect 202650 90410 202850 90480
rect 203150 90410 203350 90480
rect 203650 90410 203850 90480
rect 204150 90410 204350 90480
rect 204650 90410 204850 90480
rect 205150 90410 205350 90480
rect 205650 90410 205850 90480
rect 206150 90410 206350 90480
rect 206650 90410 206850 90480
rect 207150 90410 207350 90480
rect 207650 90410 207850 90480
rect 196020 90150 196090 90350
rect 196410 90150 196480 90350
rect 196520 90150 196590 90350
rect 196910 90150 196980 90350
rect 197020 90150 197090 90350
rect 197410 90150 197480 90350
rect 197520 90150 197590 90350
rect 197910 90150 197980 90350
rect 198020 90150 198090 90350
rect 198410 90150 198480 90350
rect 198520 90150 198590 90350
rect 198910 90150 198980 90350
rect 199020 90150 199090 90350
rect 199410 90150 199480 90350
rect 199520 90150 199590 90350
rect 199910 90150 199980 90350
rect 200020 90150 200090 90350
rect 200410 90150 200480 90350
rect 200520 90150 200590 90350
rect 200910 90150 200980 90350
rect 201020 90150 201090 90350
rect 201410 90150 201480 90350
rect 201520 90150 201590 90350
rect 201910 90150 201980 90350
rect 202020 90150 202090 90350
rect 202410 90150 202480 90350
rect 202520 90150 202590 90350
rect 202910 90150 202980 90350
rect 203020 90150 203090 90350
rect 203410 90150 203480 90350
rect 203520 90150 203590 90350
rect 203910 90150 203980 90350
rect 204020 90150 204090 90350
rect 204410 90150 204480 90350
rect 204520 90150 204590 90350
rect 204910 90150 204980 90350
rect 205020 90150 205090 90350
rect 205410 90150 205480 90350
rect 205520 90150 205590 90350
rect 205910 90150 205980 90350
rect 206020 90150 206090 90350
rect 206410 90150 206480 90350
rect 206520 90150 206590 90350
rect 206910 90150 206980 90350
rect 207020 90150 207090 90350
rect 207410 90150 207480 90350
rect 207520 90150 207590 90350
rect 207910 90150 207980 90350
rect 196150 90020 196350 90090
rect 196650 90020 196850 90090
rect 197150 90020 197350 90090
rect 197650 90020 197850 90090
rect 198150 90020 198350 90090
rect 198650 90020 198850 90090
rect 199150 90020 199350 90090
rect 199650 90020 199850 90090
rect 200150 90020 200350 90090
rect 200650 90020 200850 90090
rect 201150 90020 201350 90090
rect 201650 90020 201850 90090
rect 202150 90020 202350 90090
rect 202650 90020 202850 90090
rect 203150 90020 203350 90090
rect 203650 90020 203850 90090
rect 204150 90020 204350 90090
rect 204650 90020 204850 90090
rect 205150 90020 205350 90090
rect 205650 90020 205850 90090
rect 206150 90020 206350 90090
rect 206650 90020 206850 90090
rect 207150 90020 207350 90090
rect 207650 90020 207850 90090
rect 196150 89910 196350 89980
rect 196650 89910 196850 89980
rect 197150 89910 197350 89980
rect 197650 89910 197850 89980
rect 198150 89910 198350 89980
rect 198650 89910 198850 89980
rect 199150 89910 199350 89980
rect 199650 89910 199850 89980
rect 200150 89910 200350 89980
rect 200650 89910 200850 89980
rect 201150 89910 201350 89980
rect 201650 89910 201850 89980
rect 202150 89910 202350 89980
rect 202650 89910 202850 89980
rect 203150 89910 203350 89980
rect 203650 89910 203850 89980
rect 204150 89910 204350 89980
rect 204650 89910 204850 89980
rect 205150 89910 205350 89980
rect 205650 89910 205850 89980
rect 206150 89910 206350 89980
rect 206650 89910 206850 89980
rect 207150 89910 207350 89980
rect 207650 89910 207850 89980
rect 196020 89650 196090 89850
rect 196410 89650 196480 89850
rect 196520 89650 196590 89850
rect 196910 89650 196980 89850
rect 197020 89650 197090 89850
rect 197410 89650 197480 89850
rect 197520 89650 197590 89850
rect 197910 89650 197980 89850
rect 198020 89650 198090 89850
rect 198410 89650 198480 89850
rect 198520 89650 198590 89850
rect 198910 89650 198980 89850
rect 199020 89650 199090 89850
rect 199410 89650 199480 89850
rect 199520 89650 199590 89850
rect 199910 89650 199980 89850
rect 200020 89650 200090 89850
rect 200410 89650 200480 89850
rect 200520 89650 200590 89850
rect 200910 89650 200980 89850
rect 201020 89650 201090 89850
rect 201410 89650 201480 89850
rect 201520 89650 201590 89850
rect 201910 89650 201980 89850
rect 202020 89650 202090 89850
rect 202410 89650 202480 89850
rect 202520 89650 202590 89850
rect 202910 89650 202980 89850
rect 203020 89650 203090 89850
rect 203410 89650 203480 89850
rect 203520 89650 203590 89850
rect 203910 89650 203980 89850
rect 204020 89650 204090 89850
rect 204410 89650 204480 89850
rect 204520 89650 204590 89850
rect 204910 89650 204980 89850
rect 205020 89650 205090 89850
rect 205410 89650 205480 89850
rect 205520 89650 205590 89850
rect 205910 89650 205980 89850
rect 206020 89650 206090 89850
rect 206410 89650 206480 89850
rect 206520 89650 206590 89850
rect 206910 89650 206980 89850
rect 207020 89650 207090 89850
rect 207410 89650 207480 89850
rect 207520 89650 207590 89850
rect 207910 89650 207980 89850
rect 196150 89520 196350 89590
rect 196650 89520 196850 89590
rect 197150 89520 197350 89590
rect 197650 89520 197850 89590
rect 198150 89520 198350 89590
rect 198650 89520 198850 89590
rect 199150 89520 199350 89590
rect 199650 89520 199850 89590
rect 200150 89520 200350 89590
rect 200650 89520 200850 89590
rect 201150 89520 201350 89590
rect 201650 89520 201850 89590
rect 202150 89520 202350 89590
rect 202650 89520 202850 89590
rect 203150 89520 203350 89590
rect 203650 89520 203850 89590
rect 204150 89520 204350 89590
rect 204650 89520 204850 89590
rect 205150 89520 205350 89590
rect 205650 89520 205850 89590
rect 206150 89520 206350 89590
rect 206650 89520 206850 89590
rect 207150 89520 207350 89590
rect 207650 89520 207850 89590
rect 196150 89410 196350 89480
rect 196650 89410 196850 89480
rect 197150 89410 197350 89480
rect 197650 89410 197850 89480
rect 198150 89410 198350 89480
rect 198650 89410 198850 89480
rect 199150 89410 199350 89480
rect 199650 89410 199850 89480
rect 200150 89410 200350 89480
rect 200650 89410 200850 89480
rect 201150 89410 201350 89480
rect 201650 89410 201850 89480
rect 202150 89410 202350 89480
rect 202650 89410 202850 89480
rect 203150 89410 203350 89480
rect 203650 89410 203850 89480
rect 204150 89410 204350 89480
rect 204650 89410 204850 89480
rect 205150 89410 205350 89480
rect 205650 89410 205850 89480
rect 206150 89410 206350 89480
rect 206650 89410 206850 89480
rect 207150 89410 207350 89480
rect 207650 89410 207850 89480
rect 196020 89150 196090 89350
rect 196410 89150 196480 89350
rect 196520 89150 196590 89350
rect 196910 89150 196980 89350
rect 197020 89150 197090 89350
rect 197410 89150 197480 89350
rect 197520 89150 197590 89350
rect 197910 89150 197980 89350
rect 198020 89150 198090 89350
rect 198410 89150 198480 89350
rect 198520 89150 198590 89350
rect 198910 89150 198980 89350
rect 199020 89150 199090 89350
rect 199410 89150 199480 89350
rect 199520 89150 199590 89350
rect 199910 89150 199980 89350
rect 200020 89150 200090 89350
rect 200410 89150 200480 89350
rect 200520 89150 200590 89350
rect 200910 89150 200980 89350
rect 201020 89150 201090 89350
rect 201410 89150 201480 89350
rect 201520 89150 201590 89350
rect 201910 89150 201980 89350
rect 202020 89150 202090 89350
rect 202410 89150 202480 89350
rect 202520 89150 202590 89350
rect 202910 89150 202980 89350
rect 203020 89150 203090 89350
rect 203410 89150 203480 89350
rect 203520 89150 203590 89350
rect 203910 89150 203980 89350
rect 204020 89150 204090 89350
rect 204410 89150 204480 89350
rect 204520 89150 204590 89350
rect 204910 89150 204980 89350
rect 205020 89150 205090 89350
rect 205410 89150 205480 89350
rect 205520 89150 205590 89350
rect 205910 89150 205980 89350
rect 206020 89150 206090 89350
rect 206410 89150 206480 89350
rect 206520 89150 206590 89350
rect 206910 89150 206980 89350
rect 207020 89150 207090 89350
rect 207410 89150 207480 89350
rect 207520 89150 207590 89350
rect 207910 89150 207980 89350
rect 196150 89020 196350 89090
rect 196650 89020 196850 89090
rect 197150 89020 197350 89090
rect 197650 89020 197850 89090
rect 198150 89020 198350 89090
rect 198650 89020 198850 89090
rect 199150 89020 199350 89090
rect 199650 89020 199850 89090
rect 200150 89020 200350 89090
rect 200650 89020 200850 89090
rect 201150 89020 201350 89090
rect 201650 89020 201850 89090
rect 202150 89020 202350 89090
rect 202650 89020 202850 89090
rect 203150 89020 203350 89090
rect 203650 89020 203850 89090
rect 204150 89020 204350 89090
rect 204650 89020 204850 89090
rect 205150 89020 205350 89090
rect 205650 89020 205850 89090
rect 206150 89020 206350 89090
rect 206650 89020 206850 89090
rect 207150 89020 207350 89090
rect 207650 89020 207850 89090
rect 196150 88910 196350 88980
rect 196650 88910 196850 88980
rect 197150 88910 197350 88980
rect 197650 88910 197850 88980
rect 198150 88910 198350 88980
rect 198650 88910 198850 88980
rect 199150 88910 199350 88980
rect 199650 88910 199850 88980
rect 200150 88910 200350 88980
rect 200650 88910 200850 88980
rect 201150 88910 201350 88980
rect 201650 88910 201850 88980
rect 202150 88910 202350 88980
rect 202650 88910 202850 88980
rect 203150 88910 203350 88980
rect 203650 88910 203850 88980
rect 204150 88910 204350 88980
rect 204650 88910 204850 88980
rect 205150 88910 205350 88980
rect 205650 88910 205850 88980
rect 206150 88910 206350 88980
rect 206650 88910 206850 88980
rect 207150 88910 207350 88980
rect 207650 88910 207850 88980
rect 196020 88650 196090 88850
rect 196410 88650 196480 88850
rect 196520 88650 196590 88850
rect 196910 88650 196980 88850
rect 197020 88650 197090 88850
rect 197410 88650 197480 88850
rect 197520 88650 197590 88850
rect 197910 88650 197980 88850
rect 198020 88650 198090 88850
rect 198410 88650 198480 88850
rect 198520 88650 198590 88850
rect 198910 88650 198980 88850
rect 199020 88650 199090 88850
rect 199410 88650 199480 88850
rect 199520 88650 199590 88850
rect 199910 88650 199980 88850
rect 200020 88650 200090 88850
rect 200410 88650 200480 88850
rect 200520 88650 200590 88850
rect 200910 88650 200980 88850
rect 201020 88650 201090 88850
rect 201410 88650 201480 88850
rect 201520 88650 201590 88850
rect 201910 88650 201980 88850
rect 202020 88650 202090 88850
rect 202410 88650 202480 88850
rect 202520 88650 202590 88850
rect 202910 88650 202980 88850
rect 203020 88650 203090 88850
rect 203410 88650 203480 88850
rect 203520 88650 203590 88850
rect 203910 88650 203980 88850
rect 204020 88650 204090 88850
rect 204410 88650 204480 88850
rect 204520 88650 204590 88850
rect 204910 88650 204980 88850
rect 205020 88650 205090 88850
rect 205410 88650 205480 88850
rect 205520 88650 205590 88850
rect 205910 88650 205980 88850
rect 206020 88650 206090 88850
rect 206410 88650 206480 88850
rect 206520 88650 206590 88850
rect 206910 88650 206980 88850
rect 207020 88650 207090 88850
rect 207410 88650 207480 88850
rect 207520 88650 207590 88850
rect 207910 88650 207980 88850
rect 196150 88520 196350 88590
rect 196650 88520 196850 88590
rect 197150 88520 197350 88590
rect 197650 88520 197850 88590
rect 198150 88520 198350 88590
rect 198650 88520 198850 88590
rect 199150 88520 199350 88590
rect 199650 88520 199850 88590
rect 200150 88520 200350 88590
rect 200650 88520 200850 88590
rect 201150 88520 201350 88590
rect 201650 88520 201850 88590
rect 202150 88520 202350 88590
rect 202650 88520 202850 88590
rect 203150 88520 203350 88590
rect 203650 88520 203850 88590
rect 204150 88520 204350 88590
rect 204650 88520 204850 88590
rect 205150 88520 205350 88590
rect 205650 88520 205850 88590
rect 206150 88520 206350 88590
rect 206650 88520 206850 88590
rect 207150 88520 207350 88590
rect 207650 88520 207850 88590
rect 196150 88410 196350 88480
rect 196650 88410 196850 88480
rect 197150 88410 197350 88480
rect 197650 88410 197850 88480
rect 198150 88410 198350 88480
rect 198650 88410 198850 88480
rect 199150 88410 199350 88480
rect 199650 88410 199850 88480
rect 200150 88410 200350 88480
rect 200650 88410 200850 88480
rect 201150 88410 201350 88480
rect 201650 88410 201850 88480
rect 202150 88410 202350 88480
rect 202650 88410 202850 88480
rect 203150 88410 203350 88480
rect 203650 88410 203850 88480
rect 204150 88410 204350 88480
rect 204650 88410 204850 88480
rect 205150 88410 205350 88480
rect 205650 88410 205850 88480
rect 206150 88410 206350 88480
rect 206650 88410 206850 88480
rect 207150 88410 207350 88480
rect 207650 88410 207850 88480
rect 196020 88150 196090 88350
rect 196410 88150 196480 88350
rect 196520 88150 196590 88350
rect 196910 88150 196980 88350
rect 197020 88150 197090 88350
rect 197410 88150 197480 88350
rect 197520 88150 197590 88350
rect 197910 88150 197980 88350
rect 198020 88150 198090 88350
rect 198410 88150 198480 88350
rect 198520 88150 198590 88350
rect 198910 88150 198980 88350
rect 199020 88150 199090 88350
rect 199410 88150 199480 88350
rect 199520 88150 199590 88350
rect 199910 88150 199980 88350
rect 200020 88150 200090 88350
rect 200410 88150 200480 88350
rect 200520 88150 200590 88350
rect 200910 88150 200980 88350
rect 201020 88150 201090 88350
rect 201410 88150 201480 88350
rect 201520 88150 201590 88350
rect 201910 88150 201980 88350
rect 202020 88150 202090 88350
rect 202410 88150 202480 88350
rect 202520 88150 202590 88350
rect 202910 88150 202980 88350
rect 203020 88150 203090 88350
rect 203410 88150 203480 88350
rect 203520 88150 203590 88350
rect 203910 88150 203980 88350
rect 204020 88150 204090 88350
rect 204410 88150 204480 88350
rect 204520 88150 204590 88350
rect 204910 88150 204980 88350
rect 205020 88150 205090 88350
rect 205410 88150 205480 88350
rect 205520 88150 205590 88350
rect 205910 88150 205980 88350
rect 206020 88150 206090 88350
rect 206410 88150 206480 88350
rect 206520 88150 206590 88350
rect 206910 88150 206980 88350
rect 207020 88150 207090 88350
rect 207410 88150 207480 88350
rect 207520 88150 207590 88350
rect 207910 88150 207980 88350
rect 196150 88020 196350 88090
rect 196650 88020 196850 88090
rect 197150 88020 197350 88090
rect 197650 88020 197850 88090
rect 198150 88020 198350 88090
rect 198650 88020 198850 88090
rect 199150 88020 199350 88090
rect 199650 88020 199850 88090
rect 200150 88020 200350 88090
rect 200650 88020 200850 88090
rect 201150 88020 201350 88090
rect 201650 88020 201850 88090
rect 202150 88020 202350 88090
rect 202650 88020 202850 88090
rect 203150 88020 203350 88090
rect 203650 88020 203850 88090
rect 204150 88020 204350 88090
rect 204650 88020 204850 88090
rect 205150 88020 205350 88090
rect 205650 88020 205850 88090
rect 206150 88020 206350 88090
rect 206650 88020 206850 88090
rect 207150 88020 207350 88090
rect 207650 88020 207850 88090
rect 196150 87910 196350 87980
rect 196650 87910 196850 87980
rect 197150 87910 197350 87980
rect 197650 87910 197850 87980
rect 198150 87910 198350 87980
rect 198650 87910 198850 87980
rect 199150 87910 199350 87980
rect 199650 87910 199850 87980
rect 200150 87910 200350 87980
rect 200650 87910 200850 87980
rect 201150 87910 201350 87980
rect 201650 87910 201850 87980
rect 202150 87910 202350 87980
rect 202650 87910 202850 87980
rect 203150 87910 203350 87980
rect 203650 87910 203850 87980
rect 204150 87910 204350 87980
rect 204650 87910 204850 87980
rect 205150 87910 205350 87980
rect 205650 87910 205850 87980
rect 206150 87910 206350 87980
rect 206650 87910 206850 87980
rect 207150 87910 207350 87980
rect 207650 87910 207850 87980
rect 196020 87650 196090 87850
rect 196410 87650 196480 87850
rect 196520 87650 196590 87850
rect 196910 87650 196980 87850
rect 197020 87650 197090 87850
rect 197410 87650 197480 87850
rect 197520 87650 197590 87850
rect 197910 87650 197980 87850
rect 198020 87650 198090 87850
rect 198410 87650 198480 87850
rect 198520 87650 198590 87850
rect 198910 87650 198980 87850
rect 199020 87650 199090 87850
rect 199410 87650 199480 87850
rect 199520 87650 199590 87850
rect 199910 87650 199980 87850
rect 200020 87650 200090 87850
rect 200410 87650 200480 87850
rect 200520 87650 200590 87850
rect 200910 87650 200980 87850
rect 201020 87650 201090 87850
rect 201410 87650 201480 87850
rect 201520 87650 201590 87850
rect 201910 87650 201980 87850
rect 202020 87650 202090 87850
rect 202410 87650 202480 87850
rect 202520 87650 202590 87850
rect 202910 87650 202980 87850
rect 203020 87650 203090 87850
rect 203410 87650 203480 87850
rect 203520 87650 203590 87850
rect 203910 87650 203980 87850
rect 204020 87650 204090 87850
rect 204410 87650 204480 87850
rect 204520 87650 204590 87850
rect 204910 87650 204980 87850
rect 205020 87650 205090 87850
rect 205410 87650 205480 87850
rect 205520 87650 205590 87850
rect 205910 87650 205980 87850
rect 206020 87650 206090 87850
rect 206410 87650 206480 87850
rect 206520 87650 206590 87850
rect 206910 87650 206980 87850
rect 207020 87650 207090 87850
rect 207410 87650 207480 87850
rect 207520 87650 207590 87850
rect 207910 87650 207980 87850
rect 196150 87520 196350 87590
rect 196650 87520 196850 87590
rect 197150 87520 197350 87590
rect 197650 87520 197850 87590
rect 198150 87520 198350 87590
rect 198650 87520 198850 87590
rect 199150 87520 199350 87590
rect 199650 87520 199850 87590
rect 200150 87520 200350 87590
rect 200650 87520 200850 87590
rect 201150 87520 201350 87590
rect 201650 87520 201850 87590
rect 202150 87520 202350 87590
rect 202650 87520 202850 87590
rect 203150 87520 203350 87590
rect 203650 87520 203850 87590
rect 204150 87520 204350 87590
rect 204650 87520 204850 87590
rect 205150 87520 205350 87590
rect 205650 87520 205850 87590
rect 206150 87520 206350 87590
rect 206650 87520 206850 87590
rect 207150 87520 207350 87590
rect 207650 87520 207850 87590
rect 196150 87410 196350 87480
rect 196650 87410 196850 87480
rect 197150 87410 197350 87480
rect 197650 87410 197850 87480
rect 198150 87410 198350 87480
rect 198650 87410 198850 87480
rect 199150 87410 199350 87480
rect 199650 87410 199850 87480
rect 200150 87410 200350 87480
rect 200650 87410 200850 87480
rect 201150 87410 201350 87480
rect 201650 87410 201850 87480
rect 202150 87410 202350 87480
rect 202650 87410 202850 87480
rect 203150 87410 203350 87480
rect 203650 87410 203850 87480
rect 204150 87410 204350 87480
rect 204650 87410 204850 87480
rect 205150 87410 205350 87480
rect 205650 87410 205850 87480
rect 206150 87410 206350 87480
rect 206650 87410 206850 87480
rect 207150 87410 207350 87480
rect 207650 87410 207850 87480
rect 196020 87150 196090 87350
rect 196410 87150 196480 87350
rect 196520 87150 196590 87350
rect 196910 87150 196980 87350
rect 197020 87150 197090 87350
rect 197410 87150 197480 87350
rect 197520 87150 197590 87350
rect 197910 87150 197980 87350
rect 198020 87150 198090 87350
rect 198410 87150 198480 87350
rect 198520 87150 198590 87350
rect 198910 87150 198980 87350
rect 199020 87150 199090 87350
rect 199410 87150 199480 87350
rect 199520 87150 199590 87350
rect 199910 87150 199980 87350
rect 200020 87150 200090 87350
rect 200410 87150 200480 87350
rect 200520 87150 200590 87350
rect 200910 87150 200980 87350
rect 201020 87150 201090 87350
rect 201410 87150 201480 87350
rect 201520 87150 201590 87350
rect 201910 87150 201980 87350
rect 202020 87150 202090 87350
rect 202410 87150 202480 87350
rect 202520 87150 202590 87350
rect 202910 87150 202980 87350
rect 203020 87150 203090 87350
rect 203410 87150 203480 87350
rect 203520 87150 203590 87350
rect 203910 87150 203980 87350
rect 204020 87150 204090 87350
rect 204410 87150 204480 87350
rect 204520 87150 204590 87350
rect 204910 87150 204980 87350
rect 205020 87150 205090 87350
rect 205410 87150 205480 87350
rect 205520 87150 205590 87350
rect 205910 87150 205980 87350
rect 206020 87150 206090 87350
rect 206410 87150 206480 87350
rect 206520 87150 206590 87350
rect 206910 87150 206980 87350
rect 207020 87150 207090 87350
rect 207410 87150 207480 87350
rect 207520 87150 207590 87350
rect 207910 87150 207980 87350
rect 128760 86870 128900 87110
rect 129080 86870 129220 87110
rect 196150 87020 196350 87090
rect 196650 87020 196850 87090
rect 197150 87020 197350 87090
rect 197650 87020 197850 87090
rect 198150 87020 198350 87090
rect 198650 87020 198850 87090
rect 199150 87020 199350 87090
rect 199650 87020 199850 87090
rect 200150 87020 200350 87090
rect 200650 87020 200850 87090
rect 201150 87020 201350 87090
rect 201650 87020 201850 87090
rect 202150 87020 202350 87090
rect 202650 87020 202850 87090
rect 203150 87020 203350 87090
rect 203650 87020 203850 87090
rect 204150 87020 204350 87090
rect 204650 87020 204850 87090
rect 205150 87020 205350 87090
rect 205650 87020 205850 87090
rect 206150 87020 206350 87090
rect 206650 87020 206850 87090
rect 207150 87020 207350 87090
rect 207650 87020 207850 87090
rect 196150 86910 196350 86980
rect 196650 86910 196850 86980
rect 197150 86910 197350 86980
rect 197650 86910 197850 86980
rect 198150 86910 198350 86980
rect 198650 86910 198850 86980
rect 199150 86910 199350 86980
rect 199650 86910 199850 86980
rect 200150 86910 200350 86980
rect 200650 86910 200850 86980
rect 201150 86910 201350 86980
rect 201650 86910 201850 86980
rect 202150 86910 202350 86980
rect 202650 86910 202850 86980
rect 203150 86910 203350 86980
rect 203650 86910 203850 86980
rect 204150 86910 204350 86980
rect 204650 86910 204850 86980
rect 205150 86910 205350 86980
rect 205650 86910 205850 86980
rect 206150 86910 206350 86980
rect 206650 86910 206850 86980
rect 207150 86910 207350 86980
rect 207650 86910 207850 86980
rect 196020 86650 196090 86850
rect 128870 86510 129030 86630
rect 196410 86650 196480 86850
rect 196520 86650 196590 86850
rect 196910 86650 196980 86850
rect 197020 86650 197090 86850
rect 197410 86650 197480 86850
rect 197520 86650 197590 86850
rect 197910 86650 197980 86850
rect 198020 86650 198090 86850
rect 198410 86650 198480 86850
rect 198520 86650 198590 86850
rect 198910 86650 198980 86850
rect 199020 86650 199090 86850
rect 199410 86650 199480 86850
rect 199520 86650 199590 86850
rect 199910 86650 199980 86850
rect 200020 86650 200090 86850
rect 200410 86650 200480 86850
rect 200520 86650 200590 86850
rect 200910 86650 200980 86850
rect 201020 86650 201090 86850
rect 201410 86650 201480 86850
rect 201520 86650 201590 86850
rect 201910 86650 201980 86850
rect 202020 86650 202090 86850
rect 202410 86650 202480 86850
rect 202520 86650 202590 86850
rect 202910 86650 202980 86850
rect 203020 86650 203090 86850
rect 203410 86650 203480 86850
rect 203520 86650 203590 86850
rect 203910 86650 203980 86850
rect 204020 86650 204090 86850
rect 204410 86650 204480 86850
rect 204520 86650 204590 86850
rect 204910 86650 204980 86850
rect 205020 86650 205090 86850
rect 205410 86650 205480 86850
rect 205520 86650 205590 86850
rect 205910 86650 205980 86850
rect 206020 86650 206090 86850
rect 206410 86650 206480 86850
rect 206520 86650 206590 86850
rect 206910 86650 206980 86850
rect 207020 86650 207090 86850
rect 207410 86650 207480 86850
rect 207520 86650 207590 86850
rect 207910 86650 207980 86850
rect 196150 86520 196350 86590
rect 196650 86520 196850 86590
rect 197150 86520 197350 86590
rect 197650 86520 197850 86590
rect 198150 86520 198350 86590
rect 198650 86520 198850 86590
rect 199150 86520 199350 86590
rect 199650 86520 199850 86590
rect 200150 86520 200350 86590
rect 200650 86520 200850 86590
rect 201150 86520 201350 86590
rect 201650 86520 201850 86590
rect 202150 86520 202350 86590
rect 202650 86520 202850 86590
rect 203150 86520 203350 86590
rect 203650 86520 203850 86590
rect 204150 86520 204350 86590
rect 204650 86520 204850 86590
rect 205150 86520 205350 86590
rect 205650 86520 205850 86590
rect 206150 86520 206350 86590
rect 206650 86520 206850 86590
rect 207150 86520 207350 86590
rect 207650 86520 207850 86590
rect 196150 86410 196350 86480
rect 196650 86410 196850 86480
rect 197150 86410 197350 86480
rect 197650 86410 197850 86480
rect 198150 86410 198350 86480
rect 198650 86410 198850 86480
rect 199150 86410 199350 86480
rect 199650 86410 199850 86480
rect 200150 86410 200350 86480
rect 200650 86410 200850 86480
rect 201150 86410 201350 86480
rect 201650 86410 201850 86480
rect 202150 86410 202350 86480
rect 202650 86410 202850 86480
rect 203150 86410 203350 86480
rect 203650 86410 203850 86480
rect 204150 86410 204350 86480
rect 204650 86410 204850 86480
rect 205150 86410 205350 86480
rect 205650 86410 205850 86480
rect 206150 86410 206350 86480
rect 206650 86410 206850 86480
rect 207150 86410 207350 86480
rect 207650 86410 207850 86480
rect 196020 86150 196090 86350
rect 196410 86150 196480 86350
rect 196520 86150 196590 86350
rect 196910 86150 196980 86350
rect 197020 86150 197090 86350
rect 197410 86150 197480 86350
rect 197520 86150 197590 86350
rect 197910 86150 197980 86350
rect 198020 86150 198090 86350
rect 198410 86150 198480 86350
rect 198520 86150 198590 86350
rect 198910 86150 198980 86350
rect 199020 86150 199090 86350
rect 199410 86150 199480 86350
rect 199520 86150 199590 86350
rect 199910 86150 199980 86350
rect 200020 86150 200090 86350
rect 200410 86150 200480 86350
rect 200520 86150 200590 86350
rect 200910 86150 200980 86350
rect 201020 86150 201090 86350
rect 201410 86150 201480 86350
rect 201520 86150 201590 86350
rect 201910 86150 201980 86350
rect 202020 86150 202090 86350
rect 202410 86150 202480 86350
rect 202520 86150 202590 86350
rect 202910 86150 202980 86350
rect 203020 86150 203090 86350
rect 203410 86150 203480 86350
rect 203520 86150 203590 86350
rect 203910 86150 203980 86350
rect 204020 86150 204090 86350
rect 204410 86150 204480 86350
rect 204520 86150 204590 86350
rect 204910 86150 204980 86350
rect 205020 86150 205090 86350
rect 205410 86150 205480 86350
rect 205520 86150 205590 86350
rect 205910 86150 205980 86350
rect 206020 86150 206090 86350
rect 206410 86150 206480 86350
rect 206520 86150 206590 86350
rect 206910 86150 206980 86350
rect 207020 86150 207090 86350
rect 207410 86150 207480 86350
rect 207520 86150 207590 86350
rect 207910 86150 207980 86350
rect 196150 86020 196350 86090
rect 196650 86020 196850 86090
rect 197150 86020 197350 86090
rect 197650 86020 197850 86090
rect 198150 86020 198350 86090
rect 198650 86020 198850 86090
rect 199150 86020 199350 86090
rect 199650 86020 199850 86090
rect 200150 86020 200350 86090
rect 200650 86020 200850 86090
rect 201150 86020 201350 86090
rect 201650 86020 201850 86090
rect 202150 86020 202350 86090
rect 202650 86020 202850 86090
rect 203150 86020 203350 86090
rect 203650 86020 203850 86090
rect 204150 86020 204350 86090
rect 204650 86020 204850 86090
rect 205150 86020 205350 86090
rect 205650 86020 205850 86090
rect 206150 86020 206350 86090
rect 206650 86020 206850 86090
rect 207150 86020 207350 86090
rect 207650 86020 207850 86090
rect 196150 85910 196350 85980
rect 196650 85910 196850 85980
rect 197150 85910 197350 85980
rect 197650 85910 197850 85980
rect 198150 85910 198350 85980
rect 198650 85910 198850 85980
rect 199150 85910 199350 85980
rect 199650 85910 199850 85980
rect 200150 85910 200350 85980
rect 200650 85910 200850 85980
rect 201150 85910 201350 85980
rect 201650 85910 201850 85980
rect 202150 85910 202350 85980
rect 202650 85910 202850 85980
rect 203150 85910 203350 85980
rect 203650 85910 203850 85980
rect 204150 85910 204350 85980
rect 204650 85910 204850 85980
rect 205150 85910 205350 85980
rect 205650 85910 205850 85980
rect 206150 85910 206350 85980
rect 206650 85910 206850 85980
rect 207150 85910 207350 85980
rect 207650 85910 207850 85980
rect 196020 85650 196090 85850
rect 196410 85650 196480 85850
rect 196520 85650 196590 85850
rect 196910 85650 196980 85850
rect 197020 85650 197090 85850
rect 197410 85650 197480 85850
rect 197520 85650 197590 85850
rect 197910 85650 197980 85850
rect 198020 85650 198090 85850
rect 198410 85650 198480 85850
rect 198520 85650 198590 85850
rect 198910 85650 198980 85850
rect 199020 85650 199090 85850
rect 199410 85650 199480 85850
rect 199520 85650 199590 85850
rect 199910 85650 199980 85850
rect 200020 85650 200090 85850
rect 200410 85650 200480 85850
rect 200520 85650 200590 85850
rect 200910 85650 200980 85850
rect 201020 85650 201090 85850
rect 201410 85650 201480 85850
rect 201520 85650 201590 85850
rect 201910 85650 201980 85850
rect 202020 85650 202090 85850
rect 202410 85650 202480 85850
rect 202520 85650 202590 85850
rect 202910 85650 202980 85850
rect 203020 85650 203090 85850
rect 203410 85650 203480 85850
rect 203520 85650 203590 85850
rect 203910 85650 203980 85850
rect 204020 85650 204090 85850
rect 204410 85650 204480 85850
rect 204520 85650 204590 85850
rect 204910 85650 204980 85850
rect 205020 85650 205090 85850
rect 205410 85650 205480 85850
rect 205520 85650 205590 85850
rect 205910 85650 205980 85850
rect 206020 85650 206090 85850
rect 206410 85650 206480 85850
rect 206520 85650 206590 85850
rect 206910 85650 206980 85850
rect 207020 85650 207090 85850
rect 207410 85650 207480 85850
rect 207520 85650 207590 85850
rect 207910 85650 207980 85850
rect 196150 85520 196350 85590
rect 196650 85520 196850 85590
rect 197150 85520 197350 85590
rect 197650 85520 197850 85590
rect 198150 85520 198350 85590
rect 198650 85520 198850 85590
rect 199150 85520 199350 85590
rect 199650 85520 199850 85590
rect 200150 85520 200350 85590
rect 200650 85520 200850 85590
rect 201150 85520 201350 85590
rect 201650 85520 201850 85590
rect 202150 85520 202350 85590
rect 202650 85520 202850 85590
rect 203150 85520 203350 85590
rect 203650 85520 203850 85590
rect 204150 85520 204350 85590
rect 204650 85520 204850 85590
rect 205150 85520 205350 85590
rect 205650 85520 205850 85590
rect 206150 85520 206350 85590
rect 206650 85520 206850 85590
rect 207150 85520 207350 85590
rect 207650 85520 207850 85590
rect 196150 85410 196350 85480
rect 196650 85410 196850 85480
rect 197150 85410 197350 85480
rect 197650 85410 197850 85480
rect 198150 85410 198350 85480
rect 198650 85410 198850 85480
rect 199150 85410 199350 85480
rect 199650 85410 199850 85480
rect 200150 85410 200350 85480
rect 200650 85410 200850 85480
rect 201150 85410 201350 85480
rect 201650 85410 201850 85480
rect 202150 85410 202350 85480
rect 202650 85410 202850 85480
rect 203150 85410 203350 85480
rect 203650 85410 203850 85480
rect 204150 85410 204350 85480
rect 204650 85410 204850 85480
rect 205150 85410 205350 85480
rect 205650 85410 205850 85480
rect 206150 85410 206350 85480
rect 206650 85410 206850 85480
rect 207150 85410 207350 85480
rect 207650 85410 207850 85480
rect 196020 85150 196090 85350
rect 196410 85150 196480 85350
rect 196520 85150 196590 85350
rect 196910 85150 196980 85350
rect 197020 85150 197090 85350
rect 197410 85150 197480 85350
rect 197520 85150 197590 85350
rect 197910 85150 197980 85350
rect 198020 85150 198090 85350
rect 198410 85150 198480 85350
rect 198520 85150 198590 85350
rect 198910 85150 198980 85350
rect 199020 85150 199090 85350
rect 199410 85150 199480 85350
rect 199520 85150 199590 85350
rect 199910 85150 199980 85350
rect 200020 85150 200090 85350
rect 200410 85150 200480 85350
rect 200520 85150 200590 85350
rect 200910 85150 200980 85350
rect 201020 85150 201090 85350
rect 201410 85150 201480 85350
rect 201520 85150 201590 85350
rect 201910 85150 201980 85350
rect 202020 85150 202090 85350
rect 202410 85150 202480 85350
rect 202520 85150 202590 85350
rect 202910 85150 202980 85350
rect 203020 85150 203090 85350
rect 203410 85150 203480 85350
rect 203520 85150 203590 85350
rect 203910 85150 203980 85350
rect 204020 85150 204090 85350
rect 204410 85150 204480 85350
rect 204520 85150 204590 85350
rect 204910 85150 204980 85350
rect 205020 85150 205090 85350
rect 205410 85150 205480 85350
rect 205520 85150 205590 85350
rect 205910 85150 205980 85350
rect 206020 85150 206090 85350
rect 206410 85150 206480 85350
rect 206520 85150 206590 85350
rect 206910 85150 206980 85350
rect 207020 85150 207090 85350
rect 207410 85150 207480 85350
rect 207520 85150 207590 85350
rect 207910 85150 207980 85350
rect 196150 85020 196350 85090
rect 196650 85020 196850 85090
rect 197150 85020 197350 85090
rect 197650 85020 197850 85090
rect 198150 85020 198350 85090
rect 198650 85020 198850 85090
rect 199150 85020 199350 85090
rect 199650 85020 199850 85090
rect 200150 85020 200350 85090
rect 200650 85020 200850 85090
rect 201150 85020 201350 85090
rect 201650 85020 201850 85090
rect 202150 85020 202350 85090
rect 202650 85020 202850 85090
rect 203150 85020 203350 85090
rect 203650 85020 203850 85090
rect 204150 85020 204350 85090
rect 204650 85020 204850 85090
rect 205150 85020 205350 85090
rect 205650 85020 205850 85090
rect 206150 85020 206350 85090
rect 206650 85020 206850 85090
rect 207150 85020 207350 85090
rect 207650 85020 207850 85090
rect 196150 84910 196350 84980
rect 196650 84910 196850 84980
rect 197150 84910 197350 84980
rect 197650 84910 197850 84980
rect 198150 84910 198350 84980
rect 198650 84910 198850 84980
rect 199150 84910 199350 84980
rect 199650 84910 199850 84980
rect 200150 84910 200350 84980
rect 200650 84910 200850 84980
rect 201150 84910 201350 84980
rect 201650 84910 201850 84980
rect 202150 84910 202350 84980
rect 202650 84910 202850 84980
rect 203150 84910 203350 84980
rect 203650 84910 203850 84980
rect 204150 84910 204350 84980
rect 204650 84910 204850 84980
rect 205150 84910 205350 84980
rect 205650 84910 205850 84980
rect 206150 84910 206350 84980
rect 206650 84910 206850 84980
rect 207150 84910 207350 84980
rect 207650 84910 207850 84980
rect 196020 84650 196090 84850
rect 196410 84650 196480 84850
rect 196520 84650 196590 84850
rect 196910 84650 196980 84850
rect 197020 84650 197090 84850
rect 197410 84650 197480 84850
rect 197520 84650 197590 84850
rect 197910 84650 197980 84850
rect 198020 84650 198090 84850
rect 198410 84650 198480 84850
rect 198520 84650 198590 84850
rect 198910 84650 198980 84850
rect 199020 84650 199090 84850
rect 199410 84650 199480 84850
rect 199520 84650 199590 84850
rect 199910 84650 199980 84850
rect 200020 84650 200090 84850
rect 200410 84650 200480 84850
rect 200520 84650 200590 84850
rect 200910 84650 200980 84850
rect 201020 84650 201090 84850
rect 201410 84650 201480 84850
rect 201520 84650 201590 84850
rect 201910 84650 201980 84850
rect 202020 84650 202090 84850
rect 202410 84650 202480 84850
rect 202520 84650 202590 84850
rect 202910 84650 202980 84850
rect 203020 84650 203090 84850
rect 203410 84650 203480 84850
rect 203520 84650 203590 84850
rect 203910 84650 203980 84850
rect 204020 84650 204090 84850
rect 204410 84650 204480 84850
rect 204520 84650 204590 84850
rect 204910 84650 204980 84850
rect 205020 84650 205090 84850
rect 205410 84650 205480 84850
rect 205520 84650 205590 84850
rect 205910 84650 205980 84850
rect 206020 84650 206090 84850
rect 206410 84650 206480 84850
rect 206520 84650 206590 84850
rect 206910 84650 206980 84850
rect 207020 84650 207090 84850
rect 207410 84650 207480 84850
rect 207520 84650 207590 84850
rect 207910 84650 207980 84850
rect 196150 84520 196350 84590
rect 196650 84520 196850 84590
rect 197150 84520 197350 84590
rect 197650 84520 197850 84590
rect 198150 84520 198350 84590
rect 198650 84520 198850 84590
rect 199150 84520 199350 84590
rect 199650 84520 199850 84590
rect 200150 84520 200350 84590
rect 200650 84520 200850 84590
rect 201150 84520 201350 84590
rect 201650 84520 201850 84590
rect 202150 84520 202350 84590
rect 202650 84520 202850 84590
rect 203150 84520 203350 84590
rect 203650 84520 203850 84590
rect 204150 84520 204350 84590
rect 204650 84520 204850 84590
rect 205150 84520 205350 84590
rect 205650 84520 205850 84590
rect 206150 84520 206350 84590
rect 206650 84520 206850 84590
rect 207150 84520 207350 84590
rect 207650 84520 207850 84590
rect 196150 84410 196350 84480
rect 196650 84410 196850 84480
rect 197150 84410 197350 84480
rect 197650 84410 197850 84480
rect 198150 84410 198350 84480
rect 198650 84410 198850 84480
rect 199150 84410 199350 84480
rect 199650 84410 199850 84480
rect 200150 84410 200350 84480
rect 200650 84410 200850 84480
rect 201150 84410 201350 84480
rect 201650 84410 201850 84480
rect 202150 84410 202350 84480
rect 202650 84410 202850 84480
rect 203150 84410 203350 84480
rect 203650 84410 203850 84480
rect 204150 84410 204350 84480
rect 204650 84410 204850 84480
rect 205150 84410 205350 84480
rect 205650 84410 205850 84480
rect 206150 84410 206350 84480
rect 206650 84410 206850 84480
rect 207150 84410 207350 84480
rect 207650 84410 207850 84480
rect 196020 84150 196090 84350
rect 196410 84150 196480 84350
rect 196520 84150 196590 84350
rect 196910 84150 196980 84350
rect 197020 84150 197090 84350
rect 197410 84150 197480 84350
rect 197520 84150 197590 84350
rect 197910 84150 197980 84350
rect 198020 84150 198090 84350
rect 198410 84150 198480 84350
rect 198520 84150 198590 84350
rect 198910 84150 198980 84350
rect 199020 84150 199090 84350
rect 199410 84150 199480 84350
rect 199520 84150 199590 84350
rect 199910 84150 199980 84350
rect 200020 84150 200090 84350
rect 200410 84150 200480 84350
rect 200520 84150 200590 84350
rect 200910 84150 200980 84350
rect 201020 84150 201090 84350
rect 201410 84150 201480 84350
rect 201520 84150 201590 84350
rect 201910 84150 201980 84350
rect 202020 84150 202090 84350
rect 202410 84150 202480 84350
rect 202520 84150 202590 84350
rect 202910 84150 202980 84350
rect 203020 84150 203090 84350
rect 203410 84150 203480 84350
rect 203520 84150 203590 84350
rect 203910 84150 203980 84350
rect 204020 84150 204090 84350
rect 204410 84150 204480 84350
rect 204520 84150 204590 84350
rect 204910 84150 204980 84350
rect 205020 84150 205090 84350
rect 205410 84150 205480 84350
rect 205520 84150 205590 84350
rect 205910 84150 205980 84350
rect 206020 84150 206090 84350
rect 206410 84150 206480 84350
rect 206520 84150 206590 84350
rect 206910 84150 206980 84350
rect 207020 84150 207090 84350
rect 207410 84150 207480 84350
rect 207520 84150 207590 84350
rect 207910 84150 207980 84350
rect 196150 84020 196350 84090
rect 196650 84020 196850 84090
rect 197150 84020 197350 84090
rect 197650 84020 197850 84090
rect 198150 84020 198350 84090
rect 198650 84020 198850 84090
rect 199150 84020 199350 84090
rect 199650 84020 199850 84090
rect 200150 84020 200350 84090
rect 200650 84020 200850 84090
rect 201150 84020 201350 84090
rect 201650 84020 201850 84090
rect 202150 84020 202350 84090
rect 202650 84020 202850 84090
rect 203150 84020 203350 84090
rect 203650 84020 203850 84090
rect 204150 84020 204350 84090
rect 204650 84020 204850 84090
rect 205150 84020 205350 84090
rect 205650 84020 205850 84090
rect 206150 84020 206350 84090
rect 206650 84020 206850 84090
rect 207150 84020 207350 84090
rect 207650 84020 207850 84090
rect 196150 83910 196350 83980
rect 196650 83910 196850 83980
rect 197150 83910 197350 83980
rect 197650 83910 197850 83980
rect 198150 83910 198350 83980
rect 198650 83910 198850 83980
rect 199150 83910 199350 83980
rect 199650 83910 199850 83980
rect 200150 83910 200350 83980
rect 200650 83910 200850 83980
rect 201150 83910 201350 83980
rect 201650 83910 201850 83980
rect 202150 83910 202350 83980
rect 202650 83910 202850 83980
rect 203150 83910 203350 83980
rect 203650 83910 203850 83980
rect 204150 83910 204350 83980
rect 204650 83910 204850 83980
rect 205150 83910 205350 83980
rect 205650 83910 205850 83980
rect 206150 83910 206350 83980
rect 206650 83910 206850 83980
rect 207150 83910 207350 83980
rect 207650 83910 207850 83980
rect 196020 83650 196090 83850
rect 196410 83650 196480 83850
rect 196520 83650 196590 83850
rect 196910 83650 196980 83850
rect 197020 83650 197090 83850
rect 197410 83650 197480 83850
rect 197520 83650 197590 83850
rect 197910 83650 197980 83850
rect 198020 83650 198090 83850
rect 198410 83650 198480 83850
rect 198520 83650 198590 83850
rect 198910 83650 198980 83850
rect 199020 83650 199090 83850
rect 199410 83650 199480 83850
rect 199520 83650 199590 83850
rect 199910 83650 199980 83850
rect 200020 83650 200090 83850
rect 200410 83650 200480 83850
rect 200520 83650 200590 83850
rect 200910 83650 200980 83850
rect 201020 83650 201090 83850
rect 201410 83650 201480 83850
rect 201520 83650 201590 83850
rect 201910 83650 201980 83850
rect 202020 83650 202090 83850
rect 202410 83650 202480 83850
rect 202520 83650 202590 83850
rect 202910 83650 202980 83850
rect 203020 83650 203090 83850
rect 203410 83650 203480 83850
rect 203520 83650 203590 83850
rect 203910 83650 203980 83850
rect 204020 83650 204090 83850
rect 204410 83650 204480 83850
rect 204520 83650 204590 83850
rect 204910 83650 204980 83850
rect 205020 83650 205090 83850
rect 205410 83650 205480 83850
rect 205520 83650 205590 83850
rect 205910 83650 205980 83850
rect 206020 83650 206090 83850
rect 206410 83650 206480 83850
rect 206520 83650 206590 83850
rect 206910 83650 206980 83850
rect 207020 83650 207090 83850
rect 207410 83650 207480 83850
rect 207520 83650 207590 83850
rect 207910 83650 207980 83850
rect 196150 83520 196350 83590
rect 196650 83520 196850 83590
rect 197150 83520 197350 83590
rect 197650 83520 197850 83590
rect 198150 83520 198350 83590
rect 198650 83520 198850 83590
rect 199150 83520 199350 83590
rect 199650 83520 199850 83590
rect 200150 83520 200350 83590
rect 200650 83520 200850 83590
rect 201150 83520 201350 83590
rect 201650 83520 201850 83590
rect 202150 83520 202350 83590
rect 202650 83520 202850 83590
rect 203150 83520 203350 83590
rect 203650 83520 203850 83590
rect 204150 83520 204350 83590
rect 204650 83520 204850 83590
rect 205150 83520 205350 83590
rect 205650 83520 205850 83590
rect 206150 83520 206350 83590
rect 206650 83520 206850 83590
rect 207150 83520 207350 83590
rect 207650 83520 207850 83590
rect 196150 83410 196350 83480
rect 196650 83410 196850 83480
rect 197150 83410 197350 83480
rect 197650 83410 197850 83480
rect 198150 83410 198350 83480
rect 198650 83410 198850 83480
rect 199150 83410 199350 83480
rect 199650 83410 199850 83480
rect 200150 83410 200350 83480
rect 200650 83410 200850 83480
rect 201150 83410 201350 83480
rect 201650 83410 201850 83480
rect 202150 83410 202350 83480
rect 202650 83410 202850 83480
rect 203150 83410 203350 83480
rect 203650 83410 203850 83480
rect 204150 83410 204350 83480
rect 204650 83410 204850 83480
rect 205150 83410 205350 83480
rect 205650 83410 205850 83480
rect 206150 83410 206350 83480
rect 206650 83410 206850 83480
rect 207150 83410 207350 83480
rect 207650 83410 207850 83480
rect 196020 83150 196090 83350
rect 196410 83150 196480 83350
rect 196520 83150 196590 83350
rect 196910 83150 196980 83350
rect 197020 83150 197090 83350
rect 197410 83150 197480 83350
rect 197520 83150 197590 83350
rect 197910 83150 197980 83350
rect 198020 83150 198090 83350
rect 198410 83150 198480 83350
rect 198520 83150 198590 83350
rect 198910 83150 198980 83350
rect 199020 83150 199090 83350
rect 199410 83150 199480 83350
rect 199520 83150 199590 83350
rect 199910 83150 199980 83350
rect 200020 83150 200090 83350
rect 200410 83150 200480 83350
rect 200520 83150 200590 83350
rect 200910 83150 200980 83350
rect 201020 83150 201090 83350
rect 201410 83150 201480 83350
rect 201520 83150 201590 83350
rect 201910 83150 201980 83350
rect 202020 83150 202090 83350
rect 202410 83150 202480 83350
rect 202520 83150 202590 83350
rect 202910 83150 202980 83350
rect 203020 83150 203090 83350
rect 203410 83150 203480 83350
rect 203520 83150 203590 83350
rect 203910 83150 203980 83350
rect 204020 83150 204090 83350
rect 204410 83150 204480 83350
rect 204520 83150 204590 83350
rect 204910 83150 204980 83350
rect 205020 83150 205090 83350
rect 205410 83150 205480 83350
rect 205520 83150 205590 83350
rect 205910 83150 205980 83350
rect 206020 83150 206090 83350
rect 206410 83150 206480 83350
rect 206520 83150 206590 83350
rect 206910 83150 206980 83350
rect 207020 83150 207090 83350
rect 207410 83150 207480 83350
rect 207520 83150 207590 83350
rect 207910 83150 207980 83350
rect 196150 83020 196350 83090
rect 196650 83020 196850 83090
rect 197150 83020 197350 83090
rect 197650 83020 197850 83090
rect 198150 83020 198350 83090
rect 198650 83020 198850 83090
rect 199150 83020 199350 83090
rect 199650 83020 199850 83090
rect 200150 83020 200350 83090
rect 200650 83020 200850 83090
rect 201150 83020 201350 83090
rect 201650 83020 201850 83090
rect 202150 83020 202350 83090
rect 202650 83020 202850 83090
rect 203150 83020 203350 83090
rect 203650 83020 203850 83090
rect 204150 83020 204350 83090
rect 204650 83020 204850 83090
rect 205150 83020 205350 83090
rect 205650 83020 205850 83090
rect 206150 83020 206350 83090
rect 206650 83020 206850 83090
rect 207150 83020 207350 83090
rect 207650 83020 207850 83090
rect 196150 82910 196350 82980
rect 196650 82910 196850 82980
rect 197150 82910 197350 82980
rect 197650 82910 197850 82980
rect 198150 82910 198350 82980
rect 198650 82910 198850 82980
rect 199150 82910 199350 82980
rect 199650 82910 199850 82980
rect 200150 82910 200350 82980
rect 200650 82910 200850 82980
rect 201150 82910 201350 82980
rect 201650 82910 201850 82980
rect 202150 82910 202350 82980
rect 202650 82910 202850 82980
rect 203150 82910 203350 82980
rect 203650 82910 203850 82980
rect 204150 82910 204350 82980
rect 204650 82910 204850 82980
rect 205150 82910 205350 82980
rect 205650 82910 205850 82980
rect 206150 82910 206350 82980
rect 206650 82910 206850 82980
rect 207150 82910 207350 82980
rect 207650 82910 207850 82980
rect 196020 82650 196090 82850
rect 196410 82650 196480 82850
rect 196520 82650 196590 82850
rect 196910 82650 196980 82850
rect 197020 82650 197090 82850
rect 197410 82650 197480 82850
rect 197520 82650 197590 82850
rect 197910 82650 197980 82850
rect 198020 82650 198090 82850
rect 198410 82650 198480 82850
rect 198520 82650 198590 82850
rect 198910 82650 198980 82850
rect 199020 82650 199090 82850
rect 199410 82650 199480 82850
rect 199520 82650 199590 82850
rect 199910 82650 199980 82850
rect 200020 82650 200090 82850
rect 200410 82650 200480 82850
rect 200520 82650 200590 82850
rect 200910 82650 200980 82850
rect 201020 82650 201090 82850
rect 201410 82650 201480 82850
rect 201520 82650 201590 82850
rect 201910 82650 201980 82850
rect 202020 82650 202090 82850
rect 202410 82650 202480 82850
rect 202520 82650 202590 82850
rect 202910 82650 202980 82850
rect 203020 82650 203090 82850
rect 203410 82650 203480 82850
rect 203520 82650 203590 82850
rect 203910 82650 203980 82850
rect 204020 82650 204090 82850
rect 204410 82650 204480 82850
rect 204520 82650 204590 82850
rect 204910 82650 204980 82850
rect 205020 82650 205090 82850
rect 205410 82650 205480 82850
rect 205520 82650 205590 82850
rect 205910 82650 205980 82850
rect 206020 82650 206090 82850
rect 206410 82650 206480 82850
rect 206520 82650 206590 82850
rect 206910 82650 206980 82850
rect 207020 82650 207090 82850
rect 207410 82650 207480 82850
rect 207520 82650 207590 82850
rect 207910 82650 207980 82850
rect 196150 82520 196350 82590
rect 196650 82520 196850 82590
rect 197150 82520 197350 82590
rect 197650 82520 197850 82590
rect 198150 82520 198350 82590
rect 198650 82520 198850 82590
rect 199150 82520 199350 82590
rect 199650 82520 199850 82590
rect 200150 82520 200350 82590
rect 200650 82520 200850 82590
rect 201150 82520 201350 82590
rect 201650 82520 201850 82590
rect 202150 82520 202350 82590
rect 202650 82520 202850 82590
rect 203150 82520 203350 82590
rect 203650 82520 203850 82590
rect 204150 82520 204350 82590
rect 204650 82520 204850 82590
rect 205150 82520 205350 82590
rect 205650 82520 205850 82590
rect 206150 82520 206350 82590
rect 206650 82520 206850 82590
rect 207150 82520 207350 82590
rect 207650 82520 207850 82590
rect 196150 82410 196350 82480
rect 196650 82410 196850 82480
rect 197150 82410 197350 82480
rect 197650 82410 197850 82480
rect 198150 82410 198350 82480
rect 198650 82410 198850 82480
rect 199150 82410 199350 82480
rect 199650 82410 199850 82480
rect 200150 82410 200350 82480
rect 200650 82410 200850 82480
rect 201150 82410 201350 82480
rect 201650 82410 201850 82480
rect 202150 82410 202350 82480
rect 202650 82410 202850 82480
rect 203150 82410 203350 82480
rect 203650 82410 203850 82480
rect 204150 82410 204350 82480
rect 204650 82410 204850 82480
rect 205150 82410 205350 82480
rect 205650 82410 205850 82480
rect 206150 82410 206350 82480
rect 206650 82410 206850 82480
rect 207150 82410 207350 82480
rect 207650 82410 207850 82480
rect 196020 82150 196090 82350
rect 196410 82150 196480 82350
rect 196520 82150 196590 82350
rect 196910 82150 196980 82350
rect 197020 82150 197090 82350
rect 197410 82150 197480 82350
rect 197520 82150 197590 82350
rect 197910 82150 197980 82350
rect 198020 82150 198090 82350
rect 198410 82150 198480 82350
rect 198520 82150 198590 82350
rect 198910 82150 198980 82350
rect 199020 82150 199090 82350
rect 199410 82150 199480 82350
rect 199520 82150 199590 82350
rect 199910 82150 199980 82350
rect 200020 82150 200090 82350
rect 200410 82150 200480 82350
rect 200520 82150 200590 82350
rect 200910 82150 200980 82350
rect 201020 82150 201090 82350
rect 201410 82150 201480 82350
rect 201520 82150 201590 82350
rect 201910 82150 201980 82350
rect 202020 82150 202090 82350
rect 202410 82150 202480 82350
rect 202520 82150 202590 82350
rect 202910 82150 202980 82350
rect 203020 82150 203090 82350
rect 203410 82150 203480 82350
rect 203520 82150 203590 82350
rect 203910 82150 203980 82350
rect 204020 82150 204090 82350
rect 204410 82150 204480 82350
rect 204520 82150 204590 82350
rect 204910 82150 204980 82350
rect 205020 82150 205090 82350
rect 205410 82150 205480 82350
rect 205520 82150 205590 82350
rect 205910 82150 205980 82350
rect 206020 82150 206090 82350
rect 206410 82150 206480 82350
rect 206520 82150 206590 82350
rect 206910 82150 206980 82350
rect 207020 82150 207090 82350
rect 207410 82150 207480 82350
rect 207520 82150 207590 82350
rect 207910 82150 207980 82350
rect 196150 82020 196350 82090
rect 196650 82020 196850 82090
rect 197150 82020 197350 82090
rect 197650 82020 197850 82090
rect 198150 82020 198350 82090
rect 198650 82020 198850 82090
rect 199150 82020 199350 82090
rect 199650 82020 199850 82090
rect 200150 82020 200350 82090
rect 200650 82020 200850 82090
rect 201150 82020 201350 82090
rect 201650 82020 201850 82090
rect 202150 82020 202350 82090
rect 202650 82020 202850 82090
rect 203150 82020 203350 82090
rect 203650 82020 203850 82090
rect 204150 82020 204350 82090
rect 204650 82020 204850 82090
rect 205150 82020 205350 82090
rect 205650 82020 205850 82090
rect 206150 82020 206350 82090
rect 206650 82020 206850 82090
rect 207150 82020 207350 82090
rect 207650 82020 207850 82090
rect 196150 81910 196350 81980
rect 196650 81910 196850 81980
rect 197150 81910 197350 81980
rect 197650 81910 197850 81980
rect 198150 81910 198350 81980
rect 198650 81910 198850 81980
rect 199150 81910 199350 81980
rect 199650 81910 199850 81980
rect 200150 81910 200350 81980
rect 200650 81910 200850 81980
rect 201150 81910 201350 81980
rect 201650 81910 201850 81980
rect 202150 81910 202350 81980
rect 202650 81910 202850 81980
rect 203150 81910 203350 81980
rect 203650 81910 203850 81980
rect 204150 81910 204350 81980
rect 204650 81910 204850 81980
rect 205150 81910 205350 81980
rect 205650 81910 205850 81980
rect 206150 81910 206350 81980
rect 206650 81910 206850 81980
rect 207150 81910 207350 81980
rect 207650 81910 207850 81980
rect 196020 81650 196090 81850
rect 196410 81650 196480 81850
rect 196520 81650 196590 81850
rect 196910 81650 196980 81850
rect 197020 81650 197090 81850
rect 197410 81650 197480 81850
rect 197520 81650 197590 81850
rect 197910 81650 197980 81850
rect 198020 81650 198090 81850
rect 198410 81650 198480 81850
rect 198520 81650 198590 81850
rect 198910 81650 198980 81850
rect 199020 81650 199090 81850
rect 199410 81650 199480 81850
rect 199520 81650 199590 81850
rect 199910 81650 199980 81850
rect 200020 81650 200090 81850
rect 200410 81650 200480 81850
rect 200520 81650 200590 81850
rect 200910 81650 200980 81850
rect 201020 81650 201090 81850
rect 201410 81650 201480 81850
rect 201520 81650 201590 81850
rect 201910 81650 201980 81850
rect 202020 81650 202090 81850
rect 202410 81650 202480 81850
rect 202520 81650 202590 81850
rect 202910 81650 202980 81850
rect 203020 81650 203090 81850
rect 203410 81650 203480 81850
rect 203520 81650 203590 81850
rect 203910 81650 203980 81850
rect 204020 81650 204090 81850
rect 204410 81650 204480 81850
rect 204520 81650 204590 81850
rect 204910 81650 204980 81850
rect 205020 81650 205090 81850
rect 205410 81650 205480 81850
rect 205520 81650 205590 81850
rect 205910 81650 205980 81850
rect 206020 81650 206090 81850
rect 206410 81650 206480 81850
rect 206520 81650 206590 81850
rect 206910 81650 206980 81850
rect 207020 81650 207090 81850
rect 207410 81650 207480 81850
rect 207520 81650 207590 81850
rect 207910 81650 207980 81850
rect 196150 81520 196350 81590
rect 196650 81520 196850 81590
rect 197150 81520 197350 81590
rect 197650 81520 197850 81590
rect 198150 81520 198350 81590
rect 198650 81520 198850 81590
rect 199150 81520 199350 81590
rect 199650 81520 199850 81590
rect 200150 81520 200350 81590
rect 200650 81520 200850 81590
rect 201150 81520 201350 81590
rect 201650 81520 201850 81590
rect 202150 81520 202350 81590
rect 202650 81520 202850 81590
rect 203150 81520 203350 81590
rect 203650 81520 203850 81590
rect 204150 81520 204350 81590
rect 204650 81520 204850 81590
rect 205150 81520 205350 81590
rect 205650 81520 205850 81590
rect 206150 81520 206350 81590
rect 206650 81520 206850 81590
rect 207150 81520 207350 81590
rect 207650 81520 207850 81590
rect 196150 81410 196350 81480
rect 196650 81410 196850 81480
rect 197150 81410 197350 81480
rect 197650 81410 197850 81480
rect 198150 81410 198350 81480
rect 198650 81410 198850 81480
rect 199150 81410 199350 81480
rect 199650 81410 199850 81480
rect 200150 81410 200350 81480
rect 200650 81410 200850 81480
rect 201150 81410 201350 81480
rect 201650 81410 201850 81480
rect 202150 81410 202350 81480
rect 202650 81410 202850 81480
rect 203150 81410 203350 81480
rect 203650 81410 203850 81480
rect 204150 81410 204350 81480
rect 204650 81410 204850 81480
rect 205150 81410 205350 81480
rect 205650 81410 205850 81480
rect 206150 81410 206350 81480
rect 206650 81410 206850 81480
rect 207150 81410 207350 81480
rect 207650 81410 207850 81480
rect 196020 81150 196090 81350
rect 196410 81150 196480 81350
rect 196520 81150 196590 81350
rect 196910 81150 196980 81350
rect 197020 81150 197090 81350
rect 197410 81150 197480 81350
rect 197520 81150 197590 81350
rect 197910 81150 197980 81350
rect 198020 81150 198090 81350
rect 198410 81150 198480 81350
rect 198520 81150 198590 81350
rect 198910 81150 198980 81350
rect 199020 81150 199090 81350
rect 199410 81150 199480 81350
rect 199520 81150 199590 81350
rect 199910 81150 199980 81350
rect 200020 81150 200090 81350
rect 200410 81150 200480 81350
rect 200520 81150 200590 81350
rect 200910 81150 200980 81350
rect 201020 81150 201090 81350
rect 201410 81150 201480 81350
rect 201520 81150 201590 81350
rect 201910 81150 201980 81350
rect 202020 81150 202090 81350
rect 202410 81150 202480 81350
rect 202520 81150 202590 81350
rect 202910 81150 202980 81350
rect 203020 81150 203090 81350
rect 203410 81150 203480 81350
rect 203520 81150 203590 81350
rect 203910 81150 203980 81350
rect 204020 81150 204090 81350
rect 204410 81150 204480 81350
rect 204520 81150 204590 81350
rect 204910 81150 204980 81350
rect 205020 81150 205090 81350
rect 205410 81150 205480 81350
rect 205520 81150 205590 81350
rect 205910 81150 205980 81350
rect 206020 81150 206090 81350
rect 206410 81150 206480 81350
rect 206520 81150 206590 81350
rect 206910 81150 206980 81350
rect 207020 81150 207090 81350
rect 207410 81150 207480 81350
rect 207520 81150 207590 81350
rect 207910 81150 207980 81350
rect 196150 81020 196350 81090
rect 196650 81020 196850 81090
rect 197150 81020 197350 81090
rect 197650 81020 197850 81090
rect 198150 81020 198350 81090
rect 198650 81020 198850 81090
rect 199150 81020 199350 81090
rect 199650 81020 199850 81090
rect 200150 81020 200350 81090
rect 200650 81020 200850 81090
rect 201150 81020 201350 81090
rect 201650 81020 201850 81090
rect 202150 81020 202350 81090
rect 202650 81020 202850 81090
rect 203150 81020 203350 81090
rect 203650 81020 203850 81090
rect 204150 81020 204350 81090
rect 204650 81020 204850 81090
rect 205150 81020 205350 81090
rect 205650 81020 205850 81090
rect 206150 81020 206350 81090
rect 206650 81020 206850 81090
rect 207150 81020 207350 81090
rect 207650 81020 207850 81090
rect 196150 80910 196350 80980
rect 196650 80910 196850 80980
rect 197150 80910 197350 80980
rect 197650 80910 197850 80980
rect 198150 80910 198350 80980
rect 198650 80910 198850 80980
rect 199150 80910 199350 80980
rect 199650 80910 199850 80980
rect 200150 80910 200350 80980
rect 200650 80910 200850 80980
rect 201150 80910 201350 80980
rect 201650 80910 201850 80980
rect 202150 80910 202350 80980
rect 202650 80910 202850 80980
rect 203150 80910 203350 80980
rect 203650 80910 203850 80980
rect 204150 80910 204350 80980
rect 204650 80910 204850 80980
rect 205150 80910 205350 80980
rect 205650 80910 205850 80980
rect 206150 80910 206350 80980
rect 206650 80910 206850 80980
rect 207150 80910 207350 80980
rect 207650 80910 207850 80980
rect 196020 80650 196090 80850
rect 196410 80650 196480 80850
rect 196520 80650 196590 80850
rect 196910 80650 196980 80850
rect 197020 80650 197090 80850
rect 197410 80650 197480 80850
rect 197520 80650 197590 80850
rect 197910 80650 197980 80850
rect 198020 80650 198090 80850
rect 198410 80650 198480 80850
rect 198520 80650 198590 80850
rect 198910 80650 198980 80850
rect 199020 80650 199090 80850
rect 199410 80650 199480 80850
rect 199520 80650 199590 80850
rect 199910 80650 199980 80850
rect 200020 80650 200090 80850
rect 200410 80650 200480 80850
rect 200520 80650 200590 80850
rect 200910 80650 200980 80850
rect 201020 80650 201090 80850
rect 201410 80650 201480 80850
rect 201520 80650 201590 80850
rect 201910 80650 201980 80850
rect 202020 80650 202090 80850
rect 202410 80650 202480 80850
rect 202520 80650 202590 80850
rect 202910 80650 202980 80850
rect 203020 80650 203090 80850
rect 203410 80650 203480 80850
rect 203520 80650 203590 80850
rect 203910 80650 203980 80850
rect 204020 80650 204090 80850
rect 204410 80650 204480 80850
rect 204520 80650 204590 80850
rect 204910 80650 204980 80850
rect 205020 80650 205090 80850
rect 205410 80650 205480 80850
rect 205520 80650 205590 80850
rect 205910 80650 205980 80850
rect 206020 80650 206090 80850
rect 206410 80650 206480 80850
rect 206520 80650 206590 80850
rect 206910 80650 206980 80850
rect 207020 80650 207090 80850
rect 207410 80650 207480 80850
rect 207520 80650 207590 80850
rect 207910 80650 207980 80850
rect 196150 80520 196350 80590
rect 196650 80520 196850 80590
rect 197150 80520 197350 80590
rect 197650 80520 197850 80590
rect 198150 80520 198350 80590
rect 198650 80520 198850 80590
rect 199150 80520 199350 80590
rect 199650 80520 199850 80590
rect 200150 80520 200350 80590
rect 200650 80520 200850 80590
rect 201150 80520 201350 80590
rect 201650 80520 201850 80590
rect 202150 80520 202350 80590
rect 202650 80520 202850 80590
rect 203150 80520 203350 80590
rect 203650 80520 203850 80590
rect 204150 80520 204350 80590
rect 204650 80520 204850 80590
rect 205150 80520 205350 80590
rect 205650 80520 205850 80590
rect 206150 80520 206350 80590
rect 206650 80520 206850 80590
rect 207150 80520 207350 80590
rect 207650 80520 207850 80590
rect 196150 80410 196350 80480
rect 196650 80410 196850 80480
rect 197150 80410 197350 80480
rect 197650 80410 197850 80480
rect 198150 80410 198350 80480
rect 198650 80410 198850 80480
rect 199150 80410 199350 80480
rect 199650 80410 199850 80480
rect 200150 80410 200350 80480
rect 200650 80410 200850 80480
rect 201150 80410 201350 80480
rect 201650 80410 201850 80480
rect 202150 80410 202350 80480
rect 202650 80410 202850 80480
rect 203150 80410 203350 80480
rect 203650 80410 203850 80480
rect 204150 80410 204350 80480
rect 204650 80410 204850 80480
rect 205150 80410 205350 80480
rect 205650 80410 205850 80480
rect 206150 80410 206350 80480
rect 206650 80410 206850 80480
rect 207150 80410 207350 80480
rect 207650 80410 207850 80480
rect 196020 80150 196090 80350
rect 196410 80150 196480 80350
rect 196520 80150 196590 80350
rect 196910 80150 196980 80350
rect 197020 80150 197090 80350
rect 197410 80150 197480 80350
rect 197520 80150 197590 80350
rect 197910 80150 197980 80350
rect 198020 80150 198090 80350
rect 198410 80150 198480 80350
rect 198520 80150 198590 80350
rect 198910 80150 198980 80350
rect 199020 80150 199090 80350
rect 199410 80150 199480 80350
rect 199520 80150 199590 80350
rect 199910 80150 199980 80350
rect 200020 80150 200090 80350
rect 200410 80150 200480 80350
rect 200520 80150 200590 80350
rect 200910 80150 200980 80350
rect 201020 80150 201090 80350
rect 201410 80150 201480 80350
rect 201520 80150 201590 80350
rect 201910 80150 201980 80350
rect 202020 80150 202090 80350
rect 202410 80150 202480 80350
rect 202520 80150 202590 80350
rect 202910 80150 202980 80350
rect 203020 80150 203090 80350
rect 203410 80150 203480 80350
rect 203520 80150 203590 80350
rect 203910 80150 203980 80350
rect 204020 80150 204090 80350
rect 204410 80150 204480 80350
rect 204520 80150 204590 80350
rect 204910 80150 204980 80350
rect 205020 80150 205090 80350
rect 205410 80150 205480 80350
rect 205520 80150 205590 80350
rect 205910 80150 205980 80350
rect 206020 80150 206090 80350
rect 206410 80150 206480 80350
rect 206520 80150 206590 80350
rect 206910 80150 206980 80350
rect 207020 80150 207090 80350
rect 207410 80150 207480 80350
rect 207520 80150 207590 80350
rect 207910 80150 207980 80350
rect 196150 80020 196350 80090
rect 196650 80020 196850 80090
rect 197150 80020 197350 80090
rect 197650 80020 197850 80090
rect 198150 80020 198350 80090
rect 198650 80020 198850 80090
rect 199150 80020 199350 80090
rect 199650 80020 199850 80090
rect 200150 80020 200350 80090
rect 200650 80020 200850 80090
rect 201150 80020 201350 80090
rect 201650 80020 201850 80090
rect 202150 80020 202350 80090
rect 202650 80020 202850 80090
rect 203150 80020 203350 80090
rect 203650 80020 203850 80090
rect 204150 80020 204350 80090
rect 204650 80020 204850 80090
rect 205150 80020 205350 80090
rect 205650 80020 205850 80090
rect 206150 80020 206350 80090
rect 206650 80020 206850 80090
rect 207150 80020 207350 80090
rect 207650 80020 207850 80090
rect 196150 79910 196350 79980
rect 196650 79910 196850 79980
rect 197150 79910 197350 79980
rect 197650 79910 197850 79980
rect 198150 79910 198350 79980
rect 198650 79910 198850 79980
rect 199150 79910 199350 79980
rect 199650 79910 199850 79980
rect 200150 79910 200350 79980
rect 200650 79910 200850 79980
rect 201150 79910 201350 79980
rect 201650 79910 201850 79980
rect 202150 79910 202350 79980
rect 202650 79910 202850 79980
rect 203150 79910 203350 79980
rect 203650 79910 203850 79980
rect 204150 79910 204350 79980
rect 204650 79910 204850 79980
rect 205150 79910 205350 79980
rect 205650 79910 205850 79980
rect 206150 79910 206350 79980
rect 206650 79910 206850 79980
rect 207150 79910 207350 79980
rect 207650 79910 207850 79980
rect 196020 79650 196090 79850
rect 196410 79650 196480 79850
rect 196520 79650 196590 79850
rect 196910 79650 196980 79850
rect 197020 79650 197090 79850
rect 197410 79650 197480 79850
rect 197520 79650 197590 79850
rect 197910 79650 197980 79850
rect 198020 79650 198090 79850
rect 198410 79650 198480 79850
rect 198520 79650 198590 79850
rect 198910 79650 198980 79850
rect 199020 79650 199090 79850
rect 199410 79650 199480 79850
rect 199520 79650 199590 79850
rect 199910 79650 199980 79850
rect 200020 79650 200090 79850
rect 200410 79650 200480 79850
rect 200520 79650 200590 79850
rect 200910 79650 200980 79850
rect 201020 79650 201090 79850
rect 201410 79650 201480 79850
rect 201520 79650 201590 79850
rect 201910 79650 201980 79850
rect 202020 79650 202090 79850
rect 202410 79650 202480 79850
rect 202520 79650 202590 79850
rect 202910 79650 202980 79850
rect 203020 79650 203090 79850
rect 203410 79650 203480 79850
rect 203520 79650 203590 79850
rect 203910 79650 203980 79850
rect 204020 79650 204090 79850
rect 204410 79650 204480 79850
rect 204520 79650 204590 79850
rect 204910 79650 204980 79850
rect 205020 79650 205090 79850
rect 205410 79650 205480 79850
rect 205520 79650 205590 79850
rect 205910 79650 205980 79850
rect 206020 79650 206090 79850
rect 206410 79650 206480 79850
rect 206520 79650 206590 79850
rect 206910 79650 206980 79850
rect 207020 79650 207090 79850
rect 207410 79650 207480 79850
rect 207520 79650 207590 79850
rect 207910 79650 207980 79850
rect 196150 79520 196350 79590
rect 196650 79520 196850 79590
rect 197150 79520 197350 79590
rect 197650 79520 197850 79590
rect 198150 79520 198350 79590
rect 198650 79520 198850 79590
rect 199150 79520 199350 79590
rect 199650 79520 199850 79590
rect 200150 79520 200350 79590
rect 200650 79520 200850 79590
rect 201150 79520 201350 79590
rect 201650 79520 201850 79590
rect 202150 79520 202350 79590
rect 202650 79520 202850 79590
rect 203150 79520 203350 79590
rect 203650 79520 203850 79590
rect 204150 79520 204350 79590
rect 204650 79520 204850 79590
rect 205150 79520 205350 79590
rect 205650 79520 205850 79590
rect 206150 79520 206350 79590
rect 206650 79520 206850 79590
rect 207150 79520 207350 79590
rect 207650 79520 207850 79590
rect 196150 79410 196350 79480
rect 196650 79410 196850 79480
rect 197150 79410 197350 79480
rect 197650 79410 197850 79480
rect 198150 79410 198350 79480
rect 198650 79410 198850 79480
rect 199150 79410 199350 79480
rect 199650 79410 199850 79480
rect 200150 79410 200350 79480
rect 200650 79410 200850 79480
rect 201150 79410 201350 79480
rect 201650 79410 201850 79480
rect 202150 79410 202350 79480
rect 202650 79410 202850 79480
rect 203150 79410 203350 79480
rect 203650 79410 203850 79480
rect 204150 79410 204350 79480
rect 204650 79410 204850 79480
rect 205150 79410 205350 79480
rect 205650 79410 205850 79480
rect 206150 79410 206350 79480
rect 206650 79410 206850 79480
rect 207150 79410 207350 79480
rect 207650 79410 207850 79480
rect 196020 79150 196090 79350
rect 196410 79150 196480 79350
rect 196520 79150 196590 79350
rect 196910 79150 196980 79350
rect 197020 79150 197090 79350
rect 197410 79150 197480 79350
rect 197520 79150 197590 79350
rect 197910 79150 197980 79350
rect 198020 79150 198090 79350
rect 198410 79150 198480 79350
rect 198520 79150 198590 79350
rect 198910 79150 198980 79350
rect 199020 79150 199090 79350
rect 199410 79150 199480 79350
rect 199520 79150 199590 79350
rect 199910 79150 199980 79350
rect 200020 79150 200090 79350
rect 200410 79150 200480 79350
rect 200520 79150 200590 79350
rect 200910 79150 200980 79350
rect 201020 79150 201090 79350
rect 201410 79150 201480 79350
rect 201520 79150 201590 79350
rect 201910 79150 201980 79350
rect 202020 79150 202090 79350
rect 202410 79150 202480 79350
rect 202520 79150 202590 79350
rect 202910 79150 202980 79350
rect 203020 79150 203090 79350
rect 203410 79150 203480 79350
rect 203520 79150 203590 79350
rect 203910 79150 203980 79350
rect 204020 79150 204090 79350
rect 204410 79150 204480 79350
rect 204520 79150 204590 79350
rect 204910 79150 204980 79350
rect 205020 79150 205090 79350
rect 205410 79150 205480 79350
rect 205520 79150 205590 79350
rect 205910 79150 205980 79350
rect 206020 79150 206090 79350
rect 206410 79150 206480 79350
rect 206520 79150 206590 79350
rect 206910 79150 206980 79350
rect 207020 79150 207090 79350
rect 207410 79150 207480 79350
rect 207520 79150 207590 79350
rect 207910 79150 207980 79350
rect 196150 79020 196350 79090
rect 196650 79020 196850 79090
rect 197150 79020 197350 79090
rect 197650 79020 197850 79090
rect 198150 79020 198350 79090
rect 198650 79020 198850 79090
rect 199150 79020 199350 79090
rect 199650 79020 199850 79090
rect 200150 79020 200350 79090
rect 200650 79020 200850 79090
rect 201150 79020 201350 79090
rect 201650 79020 201850 79090
rect 202150 79020 202350 79090
rect 202650 79020 202850 79090
rect 203150 79020 203350 79090
rect 203650 79020 203850 79090
rect 204150 79020 204350 79090
rect 204650 79020 204850 79090
rect 205150 79020 205350 79090
rect 205650 79020 205850 79090
rect 206150 79020 206350 79090
rect 206650 79020 206850 79090
rect 207150 79020 207350 79090
rect 207650 79020 207850 79090
rect 196150 78910 196350 78980
rect 196650 78910 196850 78980
rect 197150 78910 197350 78980
rect 197650 78910 197850 78980
rect 198150 78910 198350 78980
rect 198650 78910 198850 78980
rect 199150 78910 199350 78980
rect 199650 78910 199850 78980
rect 200150 78910 200350 78980
rect 200650 78910 200850 78980
rect 201150 78910 201350 78980
rect 201650 78910 201850 78980
rect 202150 78910 202350 78980
rect 202650 78910 202850 78980
rect 203150 78910 203350 78980
rect 203650 78910 203850 78980
rect 204150 78910 204350 78980
rect 204650 78910 204850 78980
rect 205150 78910 205350 78980
rect 205650 78910 205850 78980
rect 206150 78910 206350 78980
rect 206650 78910 206850 78980
rect 207150 78910 207350 78980
rect 207650 78910 207850 78980
rect 196020 78650 196090 78850
rect 196410 78650 196480 78850
rect 196520 78650 196590 78850
rect 196910 78650 196980 78850
rect 197020 78650 197090 78850
rect 197410 78650 197480 78850
rect 197520 78650 197590 78850
rect 197910 78650 197980 78850
rect 198020 78650 198090 78850
rect 198410 78650 198480 78850
rect 198520 78650 198590 78850
rect 198910 78650 198980 78850
rect 199020 78650 199090 78850
rect 199410 78650 199480 78850
rect 199520 78650 199590 78850
rect 199910 78650 199980 78850
rect 200020 78650 200090 78850
rect 200410 78650 200480 78850
rect 200520 78650 200590 78850
rect 200910 78650 200980 78850
rect 201020 78650 201090 78850
rect 201410 78650 201480 78850
rect 201520 78650 201590 78850
rect 201910 78650 201980 78850
rect 202020 78650 202090 78850
rect 202410 78650 202480 78850
rect 202520 78650 202590 78850
rect 202910 78650 202980 78850
rect 203020 78650 203090 78850
rect 203410 78650 203480 78850
rect 203520 78650 203590 78850
rect 203910 78650 203980 78850
rect 204020 78650 204090 78850
rect 204410 78650 204480 78850
rect 204520 78650 204590 78850
rect 204910 78650 204980 78850
rect 205020 78650 205090 78850
rect 205410 78650 205480 78850
rect 205520 78650 205590 78850
rect 205910 78650 205980 78850
rect 206020 78650 206090 78850
rect 206410 78650 206480 78850
rect 206520 78650 206590 78850
rect 206910 78650 206980 78850
rect 207020 78650 207090 78850
rect 207410 78650 207480 78850
rect 207520 78650 207590 78850
rect 207910 78650 207980 78850
rect 196150 78520 196350 78590
rect 196650 78520 196850 78590
rect 197150 78520 197350 78590
rect 197650 78520 197850 78590
rect 198150 78520 198350 78590
rect 198650 78520 198850 78590
rect 199150 78520 199350 78590
rect 199650 78520 199850 78590
rect 200150 78520 200350 78590
rect 200650 78520 200850 78590
rect 201150 78520 201350 78590
rect 201650 78520 201850 78590
rect 202150 78520 202350 78590
rect 202650 78520 202850 78590
rect 203150 78520 203350 78590
rect 203650 78520 203850 78590
rect 204150 78520 204350 78590
rect 204650 78520 204850 78590
rect 205150 78520 205350 78590
rect 205650 78520 205850 78590
rect 206150 78520 206350 78590
rect 206650 78520 206850 78590
rect 207150 78520 207350 78590
rect 207650 78520 207850 78590
rect 196150 78410 196350 78480
rect 196650 78410 196850 78480
rect 197150 78410 197350 78480
rect 197650 78410 197850 78480
rect 198150 78410 198350 78480
rect 198650 78410 198850 78480
rect 199150 78410 199350 78480
rect 199650 78410 199850 78480
rect 200150 78410 200350 78480
rect 200650 78410 200850 78480
rect 201150 78410 201350 78480
rect 201650 78410 201850 78480
rect 202150 78410 202350 78480
rect 202650 78410 202850 78480
rect 203150 78410 203350 78480
rect 203650 78410 203850 78480
rect 204150 78410 204350 78480
rect 204650 78410 204850 78480
rect 205150 78410 205350 78480
rect 205650 78410 205850 78480
rect 206150 78410 206350 78480
rect 206650 78410 206850 78480
rect 207150 78410 207350 78480
rect 207650 78410 207850 78480
rect 196020 78150 196090 78350
rect 196410 78150 196480 78350
rect 196520 78150 196590 78350
rect 196910 78150 196980 78350
rect 197020 78150 197090 78350
rect 197410 78150 197480 78350
rect 197520 78150 197590 78350
rect 197910 78150 197980 78350
rect 198020 78150 198090 78350
rect 198410 78150 198480 78350
rect 198520 78150 198590 78350
rect 198910 78150 198980 78350
rect 199020 78150 199090 78350
rect 199410 78150 199480 78350
rect 199520 78150 199590 78350
rect 199910 78150 199980 78350
rect 200020 78150 200090 78350
rect 200410 78150 200480 78350
rect 200520 78150 200590 78350
rect 200910 78150 200980 78350
rect 201020 78150 201090 78350
rect 201410 78150 201480 78350
rect 201520 78150 201590 78350
rect 201910 78150 201980 78350
rect 202020 78150 202090 78350
rect 202410 78150 202480 78350
rect 202520 78150 202590 78350
rect 202910 78150 202980 78350
rect 203020 78150 203090 78350
rect 203410 78150 203480 78350
rect 203520 78150 203590 78350
rect 203910 78150 203980 78350
rect 204020 78150 204090 78350
rect 204410 78150 204480 78350
rect 204520 78150 204590 78350
rect 204910 78150 204980 78350
rect 205020 78150 205090 78350
rect 205410 78150 205480 78350
rect 205520 78150 205590 78350
rect 205910 78150 205980 78350
rect 206020 78150 206090 78350
rect 206410 78150 206480 78350
rect 206520 78150 206590 78350
rect 206910 78150 206980 78350
rect 207020 78150 207090 78350
rect 207410 78150 207480 78350
rect 207520 78150 207590 78350
rect 207910 78150 207980 78350
rect 196150 78020 196350 78090
rect 196650 78020 196850 78090
rect 197150 78020 197350 78090
rect 197650 78020 197850 78090
rect 198150 78020 198350 78090
rect 198650 78020 198850 78090
rect 199150 78020 199350 78090
rect 199650 78020 199850 78090
rect 200150 78020 200350 78090
rect 200650 78020 200850 78090
rect 201150 78020 201350 78090
rect 201650 78020 201850 78090
rect 202150 78020 202350 78090
rect 202650 78020 202850 78090
rect 203150 78020 203350 78090
rect 203650 78020 203850 78090
rect 204150 78020 204350 78090
rect 204650 78020 204850 78090
rect 205150 78020 205350 78090
rect 205650 78020 205850 78090
rect 206150 78020 206350 78090
rect 206650 78020 206850 78090
rect 207150 78020 207350 78090
rect 207650 78020 207850 78090
rect 196150 77910 196350 77980
rect 196650 77910 196850 77980
rect 197150 77910 197350 77980
rect 197650 77910 197850 77980
rect 198150 77910 198350 77980
rect 198650 77910 198850 77980
rect 199150 77910 199350 77980
rect 199650 77910 199850 77980
rect 200150 77910 200350 77980
rect 200650 77910 200850 77980
rect 201150 77910 201350 77980
rect 201650 77910 201850 77980
rect 202150 77910 202350 77980
rect 202650 77910 202850 77980
rect 203150 77910 203350 77980
rect 203650 77910 203850 77980
rect 204150 77910 204350 77980
rect 204650 77910 204850 77980
rect 205150 77910 205350 77980
rect 205650 77910 205850 77980
rect 206150 77910 206350 77980
rect 206650 77910 206850 77980
rect 207150 77910 207350 77980
rect 207650 77910 207850 77980
rect 196020 77650 196090 77850
rect 196410 77650 196480 77850
rect 196520 77650 196590 77850
rect 196910 77650 196980 77850
rect 197020 77650 197090 77850
rect 197410 77650 197480 77850
rect 197520 77650 197590 77850
rect 197910 77650 197980 77850
rect 198020 77650 198090 77850
rect 198410 77650 198480 77850
rect 198520 77650 198590 77850
rect 198910 77650 198980 77850
rect 199020 77650 199090 77850
rect 199410 77650 199480 77850
rect 199520 77650 199590 77850
rect 199910 77650 199980 77850
rect 200020 77650 200090 77850
rect 200410 77650 200480 77850
rect 200520 77650 200590 77850
rect 200910 77650 200980 77850
rect 201020 77650 201090 77850
rect 201410 77650 201480 77850
rect 201520 77650 201590 77850
rect 201910 77650 201980 77850
rect 202020 77650 202090 77850
rect 202410 77650 202480 77850
rect 202520 77650 202590 77850
rect 202910 77650 202980 77850
rect 203020 77650 203090 77850
rect 203410 77650 203480 77850
rect 203520 77650 203590 77850
rect 203910 77650 203980 77850
rect 204020 77650 204090 77850
rect 204410 77650 204480 77850
rect 204520 77650 204590 77850
rect 204910 77650 204980 77850
rect 205020 77650 205090 77850
rect 205410 77650 205480 77850
rect 205520 77650 205590 77850
rect 205910 77650 205980 77850
rect 206020 77650 206090 77850
rect 206410 77650 206480 77850
rect 206520 77650 206590 77850
rect 206910 77650 206980 77850
rect 207020 77650 207090 77850
rect 207410 77650 207480 77850
rect 207520 77650 207590 77850
rect 207910 77650 207980 77850
rect 196150 77520 196350 77590
rect 196650 77520 196850 77590
rect 197150 77520 197350 77590
rect 197650 77520 197850 77590
rect 198150 77520 198350 77590
rect 198650 77520 198850 77590
rect 199150 77520 199350 77590
rect 199650 77520 199850 77590
rect 200150 77520 200350 77590
rect 200650 77520 200850 77590
rect 201150 77520 201350 77590
rect 201650 77520 201850 77590
rect 202150 77520 202350 77590
rect 202650 77520 202850 77590
rect 203150 77520 203350 77590
rect 203650 77520 203850 77590
rect 204150 77520 204350 77590
rect 204650 77520 204850 77590
rect 205150 77520 205350 77590
rect 205650 77520 205850 77590
rect 206150 77520 206350 77590
rect 206650 77520 206850 77590
rect 207150 77520 207350 77590
rect 207650 77520 207850 77590
rect 196150 77410 196350 77480
rect 196650 77410 196850 77480
rect 197150 77410 197350 77480
rect 197650 77410 197850 77480
rect 198150 77410 198350 77480
rect 198650 77410 198850 77480
rect 199150 77410 199350 77480
rect 199650 77410 199850 77480
rect 200150 77410 200350 77480
rect 200650 77410 200850 77480
rect 201150 77410 201350 77480
rect 201650 77410 201850 77480
rect 202150 77410 202350 77480
rect 202650 77410 202850 77480
rect 203150 77410 203350 77480
rect 203650 77410 203850 77480
rect 204150 77410 204350 77480
rect 204650 77410 204850 77480
rect 205150 77410 205350 77480
rect 205650 77410 205850 77480
rect 206150 77410 206350 77480
rect 206650 77410 206850 77480
rect 207150 77410 207350 77480
rect 207650 77410 207850 77480
rect 196020 77150 196090 77350
rect 196410 77150 196480 77350
rect 196520 77150 196590 77350
rect 196910 77150 196980 77350
rect 197020 77150 197090 77350
rect 197410 77150 197480 77350
rect 197520 77150 197590 77350
rect 197910 77150 197980 77350
rect 198020 77150 198090 77350
rect 198410 77150 198480 77350
rect 198520 77150 198590 77350
rect 198910 77150 198980 77350
rect 199020 77150 199090 77350
rect 199410 77150 199480 77350
rect 199520 77150 199590 77350
rect 199910 77150 199980 77350
rect 200020 77150 200090 77350
rect 200410 77150 200480 77350
rect 200520 77150 200590 77350
rect 200910 77150 200980 77350
rect 201020 77150 201090 77350
rect 201410 77150 201480 77350
rect 201520 77150 201590 77350
rect 201910 77150 201980 77350
rect 202020 77150 202090 77350
rect 202410 77150 202480 77350
rect 202520 77150 202590 77350
rect 202910 77150 202980 77350
rect 203020 77150 203090 77350
rect 203410 77150 203480 77350
rect 203520 77150 203590 77350
rect 203910 77150 203980 77350
rect 204020 77150 204090 77350
rect 204410 77150 204480 77350
rect 204520 77150 204590 77350
rect 204910 77150 204980 77350
rect 205020 77150 205090 77350
rect 205410 77150 205480 77350
rect 205520 77150 205590 77350
rect 205910 77150 205980 77350
rect 206020 77150 206090 77350
rect 206410 77150 206480 77350
rect 206520 77150 206590 77350
rect 206910 77150 206980 77350
rect 207020 77150 207090 77350
rect 207410 77150 207480 77350
rect 207520 77150 207590 77350
rect 207910 77150 207980 77350
rect 196150 77020 196350 77090
rect 196650 77020 196850 77090
rect 197150 77020 197350 77090
rect 197650 77020 197850 77090
rect 198150 77020 198350 77090
rect 198650 77020 198850 77090
rect 199150 77020 199350 77090
rect 199650 77020 199850 77090
rect 200150 77020 200350 77090
rect 200650 77020 200850 77090
rect 201150 77020 201350 77090
rect 201650 77020 201850 77090
rect 202150 77020 202350 77090
rect 202650 77020 202850 77090
rect 203150 77020 203350 77090
rect 203650 77020 203850 77090
rect 204150 77020 204350 77090
rect 204650 77020 204850 77090
rect 205150 77020 205350 77090
rect 205650 77020 205850 77090
rect 206150 77020 206350 77090
rect 206650 77020 206850 77090
rect 207150 77020 207350 77090
rect 207650 77020 207850 77090
rect 196150 76910 196350 76980
rect 196650 76910 196850 76980
rect 197150 76910 197350 76980
rect 197650 76910 197850 76980
rect 198150 76910 198350 76980
rect 198650 76910 198850 76980
rect 199150 76910 199350 76980
rect 199650 76910 199850 76980
rect 200150 76910 200350 76980
rect 200650 76910 200850 76980
rect 201150 76910 201350 76980
rect 201650 76910 201850 76980
rect 202150 76910 202350 76980
rect 202650 76910 202850 76980
rect 203150 76910 203350 76980
rect 203650 76910 203850 76980
rect 204150 76910 204350 76980
rect 204650 76910 204850 76980
rect 205150 76910 205350 76980
rect 205650 76910 205850 76980
rect 206150 76910 206350 76980
rect 206650 76910 206850 76980
rect 207150 76910 207350 76980
rect 207650 76910 207850 76980
rect 196020 76650 196090 76850
rect 196410 76650 196480 76850
rect 196520 76650 196590 76850
rect 196910 76650 196980 76850
rect 197020 76650 197090 76850
rect 197410 76650 197480 76850
rect 197520 76650 197590 76850
rect 197910 76650 197980 76850
rect 198020 76650 198090 76850
rect 198410 76650 198480 76850
rect 198520 76650 198590 76850
rect 198910 76650 198980 76850
rect 199020 76650 199090 76850
rect 199410 76650 199480 76850
rect 199520 76650 199590 76850
rect 199910 76650 199980 76850
rect 200020 76650 200090 76850
rect 200410 76650 200480 76850
rect 200520 76650 200590 76850
rect 200910 76650 200980 76850
rect 201020 76650 201090 76850
rect 201410 76650 201480 76850
rect 201520 76650 201590 76850
rect 201910 76650 201980 76850
rect 202020 76650 202090 76850
rect 202410 76650 202480 76850
rect 202520 76650 202590 76850
rect 202910 76650 202980 76850
rect 203020 76650 203090 76850
rect 203410 76650 203480 76850
rect 203520 76650 203590 76850
rect 203910 76650 203980 76850
rect 204020 76650 204090 76850
rect 204410 76650 204480 76850
rect 204520 76650 204590 76850
rect 204910 76650 204980 76850
rect 205020 76650 205090 76850
rect 205410 76650 205480 76850
rect 205520 76650 205590 76850
rect 205910 76650 205980 76850
rect 206020 76650 206090 76850
rect 206410 76650 206480 76850
rect 206520 76650 206590 76850
rect 206910 76650 206980 76850
rect 207020 76650 207090 76850
rect 207410 76650 207480 76850
rect 207520 76650 207590 76850
rect 207910 76650 207980 76850
rect 196150 76520 196350 76590
rect 196650 76520 196850 76590
rect 197150 76520 197350 76590
rect 197650 76520 197850 76590
rect 198150 76520 198350 76590
rect 198650 76520 198850 76590
rect 199150 76520 199350 76590
rect 199650 76520 199850 76590
rect 200150 76520 200350 76590
rect 200650 76520 200850 76590
rect 201150 76520 201350 76590
rect 201650 76520 201850 76590
rect 202150 76520 202350 76590
rect 202650 76520 202850 76590
rect 203150 76520 203350 76590
rect 203650 76520 203850 76590
rect 204150 76520 204350 76590
rect 204650 76520 204850 76590
rect 205150 76520 205350 76590
rect 205650 76520 205850 76590
rect 206150 76520 206350 76590
rect 206650 76520 206850 76590
rect 207150 76520 207350 76590
rect 207650 76520 207850 76590
rect 196150 76410 196350 76480
rect 196650 76410 196850 76480
rect 197150 76410 197350 76480
rect 197650 76410 197850 76480
rect 198150 76410 198350 76480
rect 198650 76410 198850 76480
rect 199150 76410 199350 76480
rect 199650 76410 199850 76480
rect 200150 76410 200350 76480
rect 200650 76410 200850 76480
rect 201150 76410 201350 76480
rect 201650 76410 201850 76480
rect 202150 76410 202350 76480
rect 202650 76410 202850 76480
rect 203150 76410 203350 76480
rect 203650 76410 203850 76480
rect 204150 76410 204350 76480
rect 204650 76410 204850 76480
rect 205150 76410 205350 76480
rect 205650 76410 205850 76480
rect 206150 76410 206350 76480
rect 206650 76410 206850 76480
rect 207150 76410 207350 76480
rect 207650 76410 207850 76480
rect 196020 76150 196090 76350
rect 196410 76150 196480 76350
rect 196520 76150 196590 76350
rect 196910 76150 196980 76350
rect 197020 76150 197090 76350
rect 197410 76150 197480 76350
rect 197520 76150 197590 76350
rect 197910 76150 197980 76350
rect 198020 76150 198090 76350
rect 198410 76150 198480 76350
rect 198520 76150 198590 76350
rect 198910 76150 198980 76350
rect 199020 76150 199090 76350
rect 199410 76150 199480 76350
rect 199520 76150 199590 76350
rect 199910 76150 199980 76350
rect 200020 76150 200090 76350
rect 200410 76150 200480 76350
rect 200520 76150 200590 76350
rect 200910 76150 200980 76350
rect 201020 76150 201090 76350
rect 201410 76150 201480 76350
rect 201520 76150 201590 76350
rect 201910 76150 201980 76350
rect 202020 76150 202090 76350
rect 202410 76150 202480 76350
rect 202520 76150 202590 76350
rect 202910 76150 202980 76350
rect 203020 76150 203090 76350
rect 203410 76150 203480 76350
rect 203520 76150 203590 76350
rect 203910 76150 203980 76350
rect 204020 76150 204090 76350
rect 204410 76150 204480 76350
rect 204520 76150 204590 76350
rect 204910 76150 204980 76350
rect 205020 76150 205090 76350
rect 205410 76150 205480 76350
rect 205520 76150 205590 76350
rect 205910 76150 205980 76350
rect 206020 76150 206090 76350
rect 206410 76150 206480 76350
rect 206520 76150 206590 76350
rect 206910 76150 206980 76350
rect 207020 76150 207090 76350
rect 207410 76150 207480 76350
rect 207520 76150 207590 76350
rect 207910 76150 207980 76350
rect 196150 76020 196350 76090
rect 196650 76020 196850 76090
rect 197150 76020 197350 76090
rect 197650 76020 197850 76090
rect 198150 76020 198350 76090
rect 198650 76020 198850 76090
rect 199150 76020 199350 76090
rect 199650 76020 199850 76090
rect 200150 76020 200350 76090
rect 200650 76020 200850 76090
rect 201150 76020 201350 76090
rect 201650 76020 201850 76090
rect 202150 76020 202350 76090
rect 202650 76020 202850 76090
rect 203150 76020 203350 76090
rect 203650 76020 203850 76090
rect 204150 76020 204350 76090
rect 204650 76020 204850 76090
rect 205150 76020 205350 76090
rect 205650 76020 205850 76090
rect 206150 76020 206350 76090
rect 206650 76020 206850 76090
rect 207150 76020 207350 76090
rect 207650 76020 207850 76090
rect 196150 75910 196350 75980
rect 196650 75910 196850 75980
rect 197150 75910 197350 75980
rect 197650 75910 197850 75980
rect 198150 75910 198350 75980
rect 198650 75910 198850 75980
rect 199150 75910 199350 75980
rect 199650 75910 199850 75980
rect 200150 75910 200350 75980
rect 200650 75910 200850 75980
rect 201150 75910 201350 75980
rect 201650 75910 201850 75980
rect 202150 75910 202350 75980
rect 202650 75910 202850 75980
rect 203150 75910 203350 75980
rect 203650 75910 203850 75980
rect 204150 75910 204350 75980
rect 204650 75910 204850 75980
rect 205150 75910 205350 75980
rect 205650 75910 205850 75980
rect 206150 75910 206350 75980
rect 206650 75910 206850 75980
rect 207150 75910 207350 75980
rect 207650 75910 207850 75980
rect 196020 75650 196090 75850
rect 196410 75650 196480 75850
rect 196520 75650 196590 75850
rect 196910 75650 196980 75850
rect 197020 75650 197090 75850
rect 197410 75650 197480 75850
rect 197520 75650 197590 75850
rect 197910 75650 197980 75850
rect 198020 75650 198090 75850
rect 198410 75650 198480 75850
rect 198520 75650 198590 75850
rect 198910 75650 198980 75850
rect 199020 75650 199090 75850
rect 199410 75650 199480 75850
rect 199520 75650 199590 75850
rect 199910 75650 199980 75850
rect 200020 75650 200090 75850
rect 200410 75650 200480 75850
rect 200520 75650 200590 75850
rect 200910 75650 200980 75850
rect 201020 75650 201090 75850
rect 201410 75650 201480 75850
rect 201520 75650 201590 75850
rect 201910 75650 201980 75850
rect 202020 75650 202090 75850
rect 202410 75650 202480 75850
rect 202520 75650 202590 75850
rect 202910 75650 202980 75850
rect 203020 75650 203090 75850
rect 203410 75650 203480 75850
rect 203520 75650 203590 75850
rect 203910 75650 203980 75850
rect 204020 75650 204090 75850
rect 204410 75650 204480 75850
rect 204520 75650 204590 75850
rect 204910 75650 204980 75850
rect 205020 75650 205090 75850
rect 205410 75650 205480 75850
rect 205520 75650 205590 75850
rect 205910 75650 205980 75850
rect 206020 75650 206090 75850
rect 206410 75650 206480 75850
rect 206520 75650 206590 75850
rect 206910 75650 206980 75850
rect 207020 75650 207090 75850
rect 207410 75650 207480 75850
rect 207520 75650 207590 75850
rect 207910 75650 207980 75850
rect 196150 75520 196350 75590
rect 196650 75520 196850 75590
rect 197150 75520 197350 75590
rect 197650 75520 197850 75590
rect 198150 75520 198350 75590
rect 198650 75520 198850 75590
rect 199150 75520 199350 75590
rect 199650 75520 199850 75590
rect 200150 75520 200350 75590
rect 200650 75520 200850 75590
rect 201150 75520 201350 75590
rect 201650 75520 201850 75590
rect 202150 75520 202350 75590
rect 202650 75520 202850 75590
rect 203150 75520 203350 75590
rect 203650 75520 203850 75590
rect 204150 75520 204350 75590
rect 204650 75520 204850 75590
rect 205150 75520 205350 75590
rect 205650 75520 205850 75590
rect 206150 75520 206350 75590
rect 206650 75520 206850 75590
rect 207150 75520 207350 75590
rect 207650 75520 207850 75590
rect 196150 75410 196350 75480
rect 196650 75410 196850 75480
rect 197150 75410 197350 75480
rect 197650 75410 197850 75480
rect 198150 75410 198350 75480
rect 198650 75410 198850 75480
rect 199150 75410 199350 75480
rect 199650 75410 199850 75480
rect 200150 75410 200350 75480
rect 200650 75410 200850 75480
rect 201150 75410 201350 75480
rect 201650 75410 201850 75480
rect 202150 75410 202350 75480
rect 202650 75410 202850 75480
rect 203150 75410 203350 75480
rect 203650 75410 203850 75480
rect 204150 75410 204350 75480
rect 204650 75410 204850 75480
rect 205150 75410 205350 75480
rect 205650 75410 205850 75480
rect 206150 75410 206350 75480
rect 206650 75410 206850 75480
rect 207150 75410 207350 75480
rect 207650 75410 207850 75480
rect 196020 75150 196090 75350
rect 196410 75150 196480 75350
rect 196520 75150 196590 75350
rect 196910 75150 196980 75350
rect 197020 75150 197090 75350
rect 197410 75150 197480 75350
rect 197520 75150 197590 75350
rect 197910 75150 197980 75350
rect 198020 75150 198090 75350
rect 198410 75150 198480 75350
rect 198520 75150 198590 75350
rect 198910 75150 198980 75350
rect 199020 75150 199090 75350
rect 199410 75150 199480 75350
rect 199520 75150 199590 75350
rect 199910 75150 199980 75350
rect 200020 75150 200090 75350
rect 200410 75150 200480 75350
rect 200520 75150 200590 75350
rect 200910 75150 200980 75350
rect 201020 75150 201090 75350
rect 201410 75150 201480 75350
rect 201520 75150 201590 75350
rect 201910 75150 201980 75350
rect 202020 75150 202090 75350
rect 202410 75150 202480 75350
rect 202520 75150 202590 75350
rect 202910 75150 202980 75350
rect 203020 75150 203090 75350
rect 203410 75150 203480 75350
rect 203520 75150 203590 75350
rect 203910 75150 203980 75350
rect 204020 75150 204090 75350
rect 204410 75150 204480 75350
rect 204520 75150 204590 75350
rect 204910 75150 204980 75350
rect 205020 75150 205090 75350
rect 205410 75150 205480 75350
rect 205520 75150 205590 75350
rect 205910 75150 205980 75350
rect 206020 75150 206090 75350
rect 206410 75150 206480 75350
rect 206520 75150 206590 75350
rect 206910 75150 206980 75350
rect 207020 75150 207090 75350
rect 207410 75150 207480 75350
rect 207520 75150 207590 75350
rect 207910 75150 207980 75350
rect 196150 75020 196350 75090
rect 196650 75020 196850 75090
rect 197150 75020 197350 75090
rect 197650 75020 197850 75090
rect 198150 75020 198350 75090
rect 198650 75020 198850 75090
rect 199150 75020 199350 75090
rect 199650 75020 199850 75090
rect 200150 75020 200350 75090
rect 200650 75020 200850 75090
rect 201150 75020 201350 75090
rect 201650 75020 201850 75090
rect 202150 75020 202350 75090
rect 202650 75020 202850 75090
rect 203150 75020 203350 75090
rect 203650 75020 203850 75090
rect 204150 75020 204350 75090
rect 204650 75020 204850 75090
rect 205150 75020 205350 75090
rect 205650 75020 205850 75090
rect 206150 75020 206350 75090
rect 206650 75020 206850 75090
rect 207150 75020 207350 75090
rect 207650 75020 207850 75090
rect 196150 74910 196350 74980
rect 196650 74910 196850 74980
rect 197150 74910 197350 74980
rect 197650 74910 197850 74980
rect 198150 74910 198350 74980
rect 198650 74910 198850 74980
rect 199150 74910 199350 74980
rect 199650 74910 199850 74980
rect 200150 74910 200350 74980
rect 200650 74910 200850 74980
rect 201150 74910 201350 74980
rect 201650 74910 201850 74980
rect 202150 74910 202350 74980
rect 202650 74910 202850 74980
rect 203150 74910 203350 74980
rect 203650 74910 203850 74980
rect 204150 74910 204350 74980
rect 204650 74910 204850 74980
rect 205150 74910 205350 74980
rect 205650 74910 205850 74980
rect 206150 74910 206350 74980
rect 206650 74910 206850 74980
rect 207150 74910 207350 74980
rect 207650 74910 207850 74980
rect 196020 74650 196090 74850
rect 196410 74650 196480 74850
rect 196520 74650 196590 74850
rect 196910 74650 196980 74850
rect 197020 74650 197090 74850
rect 197410 74650 197480 74850
rect 197520 74650 197590 74850
rect 197910 74650 197980 74850
rect 198020 74650 198090 74850
rect 198410 74650 198480 74850
rect 198520 74650 198590 74850
rect 198910 74650 198980 74850
rect 199020 74650 199090 74850
rect 199410 74650 199480 74850
rect 199520 74650 199590 74850
rect 199910 74650 199980 74850
rect 200020 74650 200090 74850
rect 200410 74650 200480 74850
rect 200520 74650 200590 74850
rect 200910 74650 200980 74850
rect 201020 74650 201090 74850
rect 201410 74650 201480 74850
rect 201520 74650 201590 74850
rect 201910 74650 201980 74850
rect 202020 74650 202090 74850
rect 202410 74650 202480 74850
rect 202520 74650 202590 74850
rect 202910 74650 202980 74850
rect 203020 74650 203090 74850
rect 203410 74650 203480 74850
rect 203520 74650 203590 74850
rect 203910 74650 203980 74850
rect 204020 74650 204090 74850
rect 204410 74650 204480 74850
rect 204520 74650 204590 74850
rect 204910 74650 204980 74850
rect 205020 74650 205090 74850
rect 205410 74650 205480 74850
rect 205520 74650 205590 74850
rect 205910 74650 205980 74850
rect 206020 74650 206090 74850
rect 206410 74650 206480 74850
rect 206520 74650 206590 74850
rect 206910 74650 206980 74850
rect 207020 74650 207090 74850
rect 207410 74650 207480 74850
rect 207520 74650 207590 74850
rect 207910 74650 207980 74850
rect 196150 74520 196350 74590
rect 196650 74520 196850 74590
rect 197150 74520 197350 74590
rect 197650 74520 197850 74590
rect 198150 74520 198350 74590
rect 198650 74520 198850 74590
rect 199150 74520 199350 74590
rect 199650 74520 199850 74590
rect 200150 74520 200350 74590
rect 200650 74520 200850 74590
rect 201150 74520 201350 74590
rect 201650 74520 201850 74590
rect 202150 74520 202350 74590
rect 202650 74520 202850 74590
rect 203150 74520 203350 74590
rect 203650 74520 203850 74590
rect 204150 74520 204350 74590
rect 204650 74520 204850 74590
rect 205150 74520 205350 74590
rect 205650 74520 205850 74590
rect 206150 74520 206350 74590
rect 206650 74520 206850 74590
rect 207150 74520 207350 74590
rect 207650 74520 207850 74590
rect 196150 74410 196350 74480
rect 196650 74410 196850 74480
rect 197150 74410 197350 74480
rect 197650 74410 197850 74480
rect 198150 74410 198350 74480
rect 198650 74410 198850 74480
rect 199150 74410 199350 74480
rect 199650 74410 199850 74480
rect 200150 74410 200350 74480
rect 200650 74410 200850 74480
rect 201150 74410 201350 74480
rect 201650 74410 201850 74480
rect 202150 74410 202350 74480
rect 202650 74410 202850 74480
rect 203150 74410 203350 74480
rect 203650 74410 203850 74480
rect 204150 74410 204350 74480
rect 204650 74410 204850 74480
rect 205150 74410 205350 74480
rect 205650 74410 205850 74480
rect 206150 74410 206350 74480
rect 206650 74410 206850 74480
rect 207150 74410 207350 74480
rect 207650 74410 207850 74480
rect 196020 74150 196090 74350
rect 196410 74150 196480 74350
rect 196520 74150 196590 74350
rect 196910 74150 196980 74350
rect 197020 74150 197090 74350
rect 197410 74150 197480 74350
rect 197520 74150 197590 74350
rect 197910 74150 197980 74350
rect 198020 74150 198090 74350
rect 198410 74150 198480 74350
rect 198520 74150 198590 74350
rect 198910 74150 198980 74350
rect 199020 74150 199090 74350
rect 199410 74150 199480 74350
rect 199520 74150 199590 74350
rect 199910 74150 199980 74350
rect 200020 74150 200090 74350
rect 200410 74150 200480 74350
rect 200520 74150 200590 74350
rect 200910 74150 200980 74350
rect 201020 74150 201090 74350
rect 201410 74150 201480 74350
rect 201520 74150 201590 74350
rect 201910 74150 201980 74350
rect 202020 74150 202090 74350
rect 202410 74150 202480 74350
rect 202520 74150 202590 74350
rect 202910 74150 202980 74350
rect 203020 74150 203090 74350
rect 203410 74150 203480 74350
rect 203520 74150 203590 74350
rect 203910 74150 203980 74350
rect 204020 74150 204090 74350
rect 204410 74150 204480 74350
rect 204520 74150 204590 74350
rect 204910 74150 204980 74350
rect 205020 74150 205090 74350
rect 205410 74150 205480 74350
rect 205520 74150 205590 74350
rect 205910 74150 205980 74350
rect 206020 74150 206090 74350
rect 206410 74150 206480 74350
rect 206520 74150 206590 74350
rect 206910 74150 206980 74350
rect 207020 74150 207090 74350
rect 207410 74150 207480 74350
rect 207520 74150 207590 74350
rect 207910 74150 207980 74350
rect 196150 74020 196350 74090
rect 196650 74020 196850 74090
rect 197150 74020 197350 74090
rect 197650 74020 197850 74090
rect 198150 74020 198350 74090
rect 198650 74020 198850 74090
rect 199150 74020 199350 74090
rect 199650 74020 199850 74090
rect 200150 74020 200350 74090
rect 200650 74020 200850 74090
rect 201150 74020 201350 74090
rect 201650 74020 201850 74090
rect 202150 74020 202350 74090
rect 202650 74020 202850 74090
rect 203150 74020 203350 74090
rect 203650 74020 203850 74090
rect 204150 74020 204350 74090
rect 204650 74020 204850 74090
rect 205150 74020 205350 74090
rect 205650 74020 205850 74090
rect 206150 74020 206350 74090
rect 206650 74020 206850 74090
rect 207150 74020 207350 74090
rect 207650 74020 207850 74090
rect 196150 73910 196350 73980
rect 196650 73910 196850 73980
rect 197150 73910 197350 73980
rect 197650 73910 197850 73980
rect 198150 73910 198350 73980
rect 198650 73910 198850 73980
rect 199150 73910 199350 73980
rect 199650 73910 199850 73980
rect 200150 73910 200350 73980
rect 200650 73910 200850 73980
rect 201150 73910 201350 73980
rect 201650 73910 201850 73980
rect 202150 73910 202350 73980
rect 202650 73910 202850 73980
rect 203150 73910 203350 73980
rect 203650 73910 203850 73980
rect 204150 73910 204350 73980
rect 204650 73910 204850 73980
rect 205150 73910 205350 73980
rect 205650 73910 205850 73980
rect 206150 73910 206350 73980
rect 206650 73910 206850 73980
rect 207150 73910 207350 73980
rect 207650 73910 207850 73980
rect 196020 73650 196090 73850
rect 196410 73650 196480 73850
rect 196520 73650 196590 73850
rect 196910 73650 196980 73850
rect 197020 73650 197090 73850
rect 197410 73650 197480 73850
rect 197520 73650 197590 73850
rect 197910 73650 197980 73850
rect 198020 73650 198090 73850
rect 198410 73650 198480 73850
rect 198520 73650 198590 73850
rect 198910 73650 198980 73850
rect 199020 73650 199090 73850
rect 199410 73650 199480 73850
rect 199520 73650 199590 73850
rect 199910 73650 199980 73850
rect 200020 73650 200090 73850
rect 200410 73650 200480 73850
rect 200520 73650 200590 73850
rect 200910 73650 200980 73850
rect 201020 73650 201090 73850
rect 201410 73650 201480 73850
rect 201520 73650 201590 73850
rect 201910 73650 201980 73850
rect 202020 73650 202090 73850
rect 202410 73650 202480 73850
rect 202520 73650 202590 73850
rect 202910 73650 202980 73850
rect 203020 73650 203090 73850
rect 203410 73650 203480 73850
rect 203520 73650 203590 73850
rect 203910 73650 203980 73850
rect 204020 73650 204090 73850
rect 204410 73650 204480 73850
rect 204520 73650 204590 73850
rect 204910 73650 204980 73850
rect 205020 73650 205090 73850
rect 205410 73650 205480 73850
rect 205520 73650 205590 73850
rect 205910 73650 205980 73850
rect 206020 73650 206090 73850
rect 206410 73650 206480 73850
rect 206520 73650 206590 73850
rect 206910 73650 206980 73850
rect 207020 73650 207090 73850
rect 207410 73650 207480 73850
rect 207520 73650 207590 73850
rect 207910 73650 207980 73850
rect 196150 73520 196350 73590
rect 196650 73520 196850 73590
rect 197150 73520 197350 73590
rect 197650 73520 197850 73590
rect 198150 73520 198350 73590
rect 198650 73520 198850 73590
rect 199150 73520 199350 73590
rect 199650 73520 199850 73590
rect 200150 73520 200350 73590
rect 200650 73520 200850 73590
rect 201150 73520 201350 73590
rect 201650 73520 201850 73590
rect 202150 73520 202350 73590
rect 202650 73520 202850 73590
rect 203150 73520 203350 73590
rect 203650 73520 203850 73590
rect 204150 73520 204350 73590
rect 204650 73520 204850 73590
rect 205150 73520 205350 73590
rect 205650 73520 205850 73590
rect 206150 73520 206350 73590
rect 206650 73520 206850 73590
rect 207150 73520 207350 73590
rect 207650 73520 207850 73590
rect 196150 73410 196350 73480
rect 196650 73410 196850 73480
rect 197150 73410 197350 73480
rect 197650 73410 197850 73480
rect 198150 73410 198350 73480
rect 198650 73410 198850 73480
rect 199150 73410 199350 73480
rect 199650 73410 199850 73480
rect 200150 73410 200350 73480
rect 200650 73410 200850 73480
rect 201150 73410 201350 73480
rect 201650 73410 201850 73480
rect 202150 73410 202350 73480
rect 202650 73410 202850 73480
rect 203150 73410 203350 73480
rect 203650 73410 203850 73480
rect 204150 73410 204350 73480
rect 204650 73410 204850 73480
rect 205150 73410 205350 73480
rect 205650 73410 205850 73480
rect 206150 73410 206350 73480
rect 206650 73410 206850 73480
rect 207150 73410 207350 73480
rect 207650 73410 207850 73480
rect 196020 73150 196090 73350
rect 196410 73150 196480 73350
rect 196520 73150 196590 73350
rect 196910 73150 196980 73350
rect 197020 73150 197090 73350
rect 197410 73150 197480 73350
rect 197520 73150 197590 73350
rect 197910 73150 197980 73350
rect 198020 73150 198090 73350
rect 198410 73150 198480 73350
rect 198520 73150 198590 73350
rect 198910 73150 198980 73350
rect 199020 73150 199090 73350
rect 199410 73150 199480 73350
rect 199520 73150 199590 73350
rect 199910 73150 199980 73350
rect 200020 73150 200090 73350
rect 200410 73150 200480 73350
rect 200520 73150 200590 73350
rect 200910 73150 200980 73350
rect 201020 73150 201090 73350
rect 201410 73150 201480 73350
rect 201520 73150 201590 73350
rect 201910 73150 201980 73350
rect 202020 73150 202090 73350
rect 202410 73150 202480 73350
rect 202520 73150 202590 73350
rect 202910 73150 202980 73350
rect 203020 73150 203090 73350
rect 203410 73150 203480 73350
rect 203520 73150 203590 73350
rect 203910 73150 203980 73350
rect 204020 73150 204090 73350
rect 204410 73150 204480 73350
rect 204520 73150 204590 73350
rect 204910 73150 204980 73350
rect 205020 73150 205090 73350
rect 205410 73150 205480 73350
rect 205520 73150 205590 73350
rect 205910 73150 205980 73350
rect 206020 73150 206090 73350
rect 206410 73150 206480 73350
rect 206520 73150 206590 73350
rect 206910 73150 206980 73350
rect 207020 73150 207090 73350
rect 207410 73150 207480 73350
rect 207520 73150 207590 73350
rect 207910 73150 207980 73350
rect 196150 73020 196350 73090
rect 196650 73020 196850 73090
rect 197150 73020 197350 73090
rect 197650 73020 197850 73090
rect 198150 73020 198350 73090
rect 198650 73020 198850 73090
rect 199150 73020 199350 73090
rect 199650 73020 199850 73090
rect 200150 73020 200350 73090
rect 200650 73020 200850 73090
rect 201150 73020 201350 73090
rect 201650 73020 201850 73090
rect 202150 73020 202350 73090
rect 202650 73020 202850 73090
rect 203150 73020 203350 73090
rect 203650 73020 203850 73090
rect 204150 73020 204350 73090
rect 204650 73020 204850 73090
rect 205150 73020 205350 73090
rect 205650 73020 205850 73090
rect 206150 73020 206350 73090
rect 206650 73020 206850 73090
rect 207150 73020 207350 73090
rect 207650 73020 207850 73090
rect 196150 72910 196350 72980
rect 196650 72910 196850 72980
rect 197150 72910 197350 72980
rect 197650 72910 197850 72980
rect 198150 72910 198350 72980
rect 198650 72910 198850 72980
rect 199150 72910 199350 72980
rect 199650 72910 199850 72980
rect 200150 72910 200350 72980
rect 200650 72910 200850 72980
rect 201150 72910 201350 72980
rect 201650 72910 201850 72980
rect 202150 72910 202350 72980
rect 202650 72910 202850 72980
rect 203150 72910 203350 72980
rect 203650 72910 203850 72980
rect 204150 72910 204350 72980
rect 204650 72910 204850 72980
rect 205150 72910 205350 72980
rect 205650 72910 205850 72980
rect 206150 72910 206350 72980
rect 206650 72910 206850 72980
rect 207150 72910 207350 72980
rect 207650 72910 207850 72980
rect 196020 72650 196090 72850
rect 196410 72650 196480 72850
rect 196520 72650 196590 72850
rect 196910 72650 196980 72850
rect 197020 72650 197090 72850
rect 197410 72650 197480 72850
rect 197520 72650 197590 72850
rect 197910 72650 197980 72850
rect 198020 72650 198090 72850
rect 198410 72650 198480 72850
rect 198520 72650 198590 72850
rect 198910 72650 198980 72850
rect 199020 72650 199090 72850
rect 199410 72650 199480 72850
rect 199520 72650 199590 72850
rect 199910 72650 199980 72850
rect 200020 72650 200090 72850
rect 200410 72650 200480 72850
rect 200520 72650 200590 72850
rect 200910 72650 200980 72850
rect 201020 72650 201090 72850
rect 201410 72650 201480 72850
rect 201520 72650 201590 72850
rect 201910 72650 201980 72850
rect 202020 72650 202090 72850
rect 202410 72650 202480 72850
rect 202520 72650 202590 72850
rect 202910 72650 202980 72850
rect 203020 72650 203090 72850
rect 203410 72650 203480 72850
rect 203520 72650 203590 72850
rect 203910 72650 203980 72850
rect 204020 72650 204090 72850
rect 204410 72650 204480 72850
rect 204520 72650 204590 72850
rect 204910 72650 204980 72850
rect 205020 72650 205090 72850
rect 205410 72650 205480 72850
rect 205520 72650 205590 72850
rect 205910 72650 205980 72850
rect 206020 72650 206090 72850
rect 206410 72650 206480 72850
rect 206520 72650 206590 72850
rect 206910 72650 206980 72850
rect 207020 72650 207090 72850
rect 207410 72650 207480 72850
rect 207520 72650 207590 72850
rect 207910 72650 207980 72850
rect 196150 72520 196350 72590
rect 196650 72520 196850 72590
rect 197150 72520 197350 72590
rect 197650 72520 197850 72590
rect 198150 72520 198350 72590
rect 198650 72520 198850 72590
rect 199150 72520 199350 72590
rect 199650 72520 199850 72590
rect 200150 72520 200350 72590
rect 200650 72520 200850 72590
rect 201150 72520 201350 72590
rect 201650 72520 201850 72590
rect 202150 72520 202350 72590
rect 202650 72520 202850 72590
rect 203150 72520 203350 72590
rect 203650 72520 203850 72590
rect 204150 72520 204350 72590
rect 204650 72520 204850 72590
rect 205150 72520 205350 72590
rect 205650 72520 205850 72590
rect 206150 72520 206350 72590
rect 206650 72520 206850 72590
rect 207150 72520 207350 72590
rect 207650 72520 207850 72590
rect 196150 72410 196350 72480
rect 196650 72410 196850 72480
rect 197150 72410 197350 72480
rect 197650 72410 197850 72480
rect 198150 72410 198350 72480
rect 198650 72410 198850 72480
rect 199150 72410 199350 72480
rect 199650 72410 199850 72480
rect 200150 72410 200350 72480
rect 200650 72410 200850 72480
rect 201150 72410 201350 72480
rect 201650 72410 201850 72480
rect 202150 72410 202350 72480
rect 202650 72410 202850 72480
rect 203150 72410 203350 72480
rect 203650 72410 203850 72480
rect 204150 72410 204350 72480
rect 204650 72410 204850 72480
rect 205150 72410 205350 72480
rect 205650 72410 205850 72480
rect 206150 72410 206350 72480
rect 206650 72410 206850 72480
rect 207150 72410 207350 72480
rect 207650 72410 207850 72480
rect 196020 72150 196090 72350
rect 196410 72150 196480 72350
rect 196520 72150 196590 72350
rect 196910 72150 196980 72350
rect 197020 72150 197090 72350
rect 197410 72150 197480 72350
rect 197520 72150 197590 72350
rect 197910 72150 197980 72350
rect 198020 72150 198090 72350
rect 198410 72150 198480 72350
rect 198520 72150 198590 72350
rect 198910 72150 198980 72350
rect 199020 72150 199090 72350
rect 199410 72150 199480 72350
rect 199520 72150 199590 72350
rect 199910 72150 199980 72350
rect 200020 72150 200090 72350
rect 200410 72150 200480 72350
rect 200520 72150 200590 72350
rect 200910 72150 200980 72350
rect 201020 72150 201090 72350
rect 201410 72150 201480 72350
rect 201520 72150 201590 72350
rect 201910 72150 201980 72350
rect 202020 72150 202090 72350
rect 202410 72150 202480 72350
rect 202520 72150 202590 72350
rect 202910 72150 202980 72350
rect 203020 72150 203090 72350
rect 203410 72150 203480 72350
rect 203520 72150 203590 72350
rect 203910 72150 203980 72350
rect 204020 72150 204090 72350
rect 204410 72150 204480 72350
rect 204520 72150 204590 72350
rect 204910 72150 204980 72350
rect 205020 72150 205090 72350
rect 205410 72150 205480 72350
rect 205520 72150 205590 72350
rect 205910 72150 205980 72350
rect 206020 72150 206090 72350
rect 206410 72150 206480 72350
rect 206520 72150 206590 72350
rect 206910 72150 206980 72350
rect 207020 72150 207090 72350
rect 207410 72150 207480 72350
rect 207520 72150 207590 72350
rect 207910 72150 207980 72350
rect 196150 72020 196350 72090
rect 196650 72020 196850 72090
rect 197150 72020 197350 72090
rect 197650 72020 197850 72090
rect 198150 72020 198350 72090
rect 198650 72020 198850 72090
rect 199150 72020 199350 72090
rect 199650 72020 199850 72090
rect 200150 72020 200350 72090
rect 200650 72020 200850 72090
rect 201150 72020 201350 72090
rect 201650 72020 201850 72090
rect 202150 72020 202350 72090
rect 202650 72020 202850 72090
rect 203150 72020 203350 72090
rect 203650 72020 203850 72090
rect 204150 72020 204350 72090
rect 204650 72020 204850 72090
rect 205150 72020 205350 72090
rect 205650 72020 205850 72090
rect 206150 72020 206350 72090
rect 206650 72020 206850 72090
rect 207150 72020 207350 72090
rect 207650 72020 207850 72090
rect 196150 71910 196350 71980
rect 196650 71910 196850 71980
rect 197150 71910 197350 71980
rect 197650 71910 197850 71980
rect 198150 71910 198350 71980
rect 198650 71910 198850 71980
rect 199150 71910 199350 71980
rect 199650 71910 199850 71980
rect 200150 71910 200350 71980
rect 200650 71910 200850 71980
rect 201150 71910 201350 71980
rect 201650 71910 201850 71980
rect 202150 71910 202350 71980
rect 202650 71910 202850 71980
rect 203150 71910 203350 71980
rect 203650 71910 203850 71980
rect 204150 71910 204350 71980
rect 204650 71910 204850 71980
rect 205150 71910 205350 71980
rect 205650 71910 205850 71980
rect 206150 71910 206350 71980
rect 206650 71910 206850 71980
rect 207150 71910 207350 71980
rect 207650 71910 207850 71980
rect 196020 71650 196090 71850
rect 196410 71650 196480 71850
rect 196520 71650 196590 71850
rect 196910 71650 196980 71850
rect 197020 71650 197090 71850
rect 197410 71650 197480 71850
rect 197520 71650 197590 71850
rect 197910 71650 197980 71850
rect 198020 71650 198090 71850
rect 198410 71650 198480 71850
rect 198520 71650 198590 71850
rect 198910 71650 198980 71850
rect 199020 71650 199090 71850
rect 199410 71650 199480 71850
rect 199520 71650 199590 71850
rect 199910 71650 199980 71850
rect 200020 71650 200090 71850
rect 200410 71650 200480 71850
rect 200520 71650 200590 71850
rect 200910 71650 200980 71850
rect 201020 71650 201090 71850
rect 201410 71650 201480 71850
rect 201520 71650 201590 71850
rect 201910 71650 201980 71850
rect 202020 71650 202090 71850
rect 202410 71650 202480 71850
rect 202520 71650 202590 71850
rect 202910 71650 202980 71850
rect 203020 71650 203090 71850
rect 203410 71650 203480 71850
rect 203520 71650 203590 71850
rect 203910 71650 203980 71850
rect 204020 71650 204090 71850
rect 204410 71650 204480 71850
rect 204520 71650 204590 71850
rect 204910 71650 204980 71850
rect 205020 71650 205090 71850
rect 205410 71650 205480 71850
rect 205520 71650 205590 71850
rect 205910 71650 205980 71850
rect 206020 71650 206090 71850
rect 206410 71650 206480 71850
rect 206520 71650 206590 71850
rect 206910 71650 206980 71850
rect 207020 71650 207090 71850
rect 207410 71650 207480 71850
rect 207520 71650 207590 71850
rect 207910 71650 207980 71850
rect 196150 71520 196350 71590
rect 196650 71520 196850 71590
rect 197150 71520 197350 71590
rect 197650 71520 197850 71590
rect 198150 71520 198350 71590
rect 198650 71520 198850 71590
rect 199150 71520 199350 71590
rect 199650 71520 199850 71590
rect 200150 71520 200350 71590
rect 200650 71520 200850 71590
rect 201150 71520 201350 71590
rect 201650 71520 201850 71590
rect 202150 71520 202350 71590
rect 202650 71520 202850 71590
rect 203150 71520 203350 71590
rect 203650 71520 203850 71590
rect 204150 71520 204350 71590
rect 204650 71520 204850 71590
rect 205150 71520 205350 71590
rect 205650 71520 205850 71590
rect 206150 71520 206350 71590
rect 206650 71520 206850 71590
rect 207150 71520 207350 71590
rect 207650 71520 207850 71590
rect 196150 71410 196350 71480
rect 196650 71410 196850 71480
rect 197150 71410 197350 71480
rect 197650 71410 197850 71480
rect 198150 71410 198350 71480
rect 198650 71410 198850 71480
rect 199150 71410 199350 71480
rect 199650 71410 199850 71480
rect 200150 71410 200350 71480
rect 200650 71410 200850 71480
rect 201150 71410 201350 71480
rect 201650 71410 201850 71480
rect 202150 71410 202350 71480
rect 202650 71410 202850 71480
rect 203150 71410 203350 71480
rect 203650 71410 203850 71480
rect 204150 71410 204350 71480
rect 204650 71410 204850 71480
rect 205150 71410 205350 71480
rect 205650 71410 205850 71480
rect 206150 71410 206350 71480
rect 206650 71410 206850 71480
rect 207150 71410 207350 71480
rect 207650 71410 207850 71480
rect 196020 71150 196090 71350
rect 196410 71150 196480 71350
rect 196520 71150 196590 71350
rect 196910 71150 196980 71350
rect 197020 71150 197090 71350
rect 197410 71150 197480 71350
rect 197520 71150 197590 71350
rect 197910 71150 197980 71350
rect 198020 71150 198090 71350
rect 198410 71150 198480 71350
rect 198520 71150 198590 71350
rect 198910 71150 198980 71350
rect 199020 71150 199090 71350
rect 199410 71150 199480 71350
rect 199520 71150 199590 71350
rect 199910 71150 199980 71350
rect 200020 71150 200090 71350
rect 200410 71150 200480 71350
rect 200520 71150 200590 71350
rect 200910 71150 200980 71350
rect 201020 71150 201090 71350
rect 201410 71150 201480 71350
rect 201520 71150 201590 71350
rect 201910 71150 201980 71350
rect 202020 71150 202090 71350
rect 202410 71150 202480 71350
rect 202520 71150 202590 71350
rect 202910 71150 202980 71350
rect 203020 71150 203090 71350
rect 203410 71150 203480 71350
rect 203520 71150 203590 71350
rect 203910 71150 203980 71350
rect 204020 71150 204090 71350
rect 204410 71150 204480 71350
rect 204520 71150 204590 71350
rect 204910 71150 204980 71350
rect 205020 71150 205090 71350
rect 205410 71150 205480 71350
rect 205520 71150 205590 71350
rect 205910 71150 205980 71350
rect 206020 71150 206090 71350
rect 206410 71150 206480 71350
rect 206520 71150 206590 71350
rect 206910 71150 206980 71350
rect 207020 71150 207090 71350
rect 207410 71150 207480 71350
rect 207520 71150 207590 71350
rect 207910 71150 207980 71350
rect 196150 71020 196350 71090
rect 196650 71020 196850 71090
rect 197150 71020 197350 71090
rect 197650 71020 197850 71090
rect 198150 71020 198350 71090
rect 198650 71020 198850 71090
rect 199150 71020 199350 71090
rect 199650 71020 199850 71090
rect 200150 71020 200350 71090
rect 200650 71020 200850 71090
rect 201150 71020 201350 71090
rect 201650 71020 201850 71090
rect 202150 71020 202350 71090
rect 202650 71020 202850 71090
rect 203150 71020 203350 71090
rect 203650 71020 203850 71090
rect 204150 71020 204350 71090
rect 204650 71020 204850 71090
rect 205150 71020 205350 71090
rect 205650 71020 205850 71090
rect 206150 71020 206350 71090
rect 206650 71020 206850 71090
rect 207150 71020 207350 71090
rect 207650 71020 207850 71090
rect 196150 70910 196350 70980
rect 196650 70910 196850 70980
rect 197150 70910 197350 70980
rect 197650 70910 197850 70980
rect 198150 70910 198350 70980
rect 198650 70910 198850 70980
rect 199150 70910 199350 70980
rect 199650 70910 199850 70980
rect 200150 70910 200350 70980
rect 200650 70910 200850 70980
rect 201150 70910 201350 70980
rect 201650 70910 201850 70980
rect 202150 70910 202350 70980
rect 202650 70910 202850 70980
rect 203150 70910 203350 70980
rect 203650 70910 203850 70980
rect 204150 70910 204350 70980
rect 204650 70910 204850 70980
rect 205150 70910 205350 70980
rect 205650 70910 205850 70980
rect 206150 70910 206350 70980
rect 206650 70910 206850 70980
rect 207150 70910 207350 70980
rect 207650 70910 207850 70980
rect 196020 70650 196090 70850
rect 196410 70650 196480 70850
rect 196520 70650 196590 70850
rect 196910 70650 196980 70850
rect 197020 70650 197090 70850
rect 197410 70650 197480 70850
rect 197520 70650 197590 70850
rect 197910 70650 197980 70850
rect 198020 70650 198090 70850
rect 198410 70650 198480 70850
rect 198520 70650 198590 70850
rect 198910 70650 198980 70850
rect 199020 70650 199090 70850
rect 199410 70650 199480 70850
rect 199520 70650 199590 70850
rect 199910 70650 199980 70850
rect 200020 70650 200090 70850
rect 200410 70650 200480 70850
rect 200520 70650 200590 70850
rect 200910 70650 200980 70850
rect 201020 70650 201090 70850
rect 201410 70650 201480 70850
rect 201520 70650 201590 70850
rect 201910 70650 201980 70850
rect 202020 70650 202090 70850
rect 202410 70650 202480 70850
rect 202520 70650 202590 70850
rect 202910 70650 202980 70850
rect 203020 70650 203090 70850
rect 203410 70650 203480 70850
rect 203520 70650 203590 70850
rect 203910 70650 203980 70850
rect 204020 70650 204090 70850
rect 204410 70650 204480 70850
rect 204520 70650 204590 70850
rect 204910 70650 204980 70850
rect 205020 70650 205090 70850
rect 205410 70650 205480 70850
rect 205520 70650 205590 70850
rect 205910 70650 205980 70850
rect 206020 70650 206090 70850
rect 206410 70650 206480 70850
rect 206520 70650 206590 70850
rect 206910 70650 206980 70850
rect 207020 70650 207090 70850
rect 207410 70650 207480 70850
rect 207520 70650 207590 70850
rect 207910 70650 207980 70850
rect 196150 70520 196350 70590
rect 196650 70520 196850 70590
rect 197150 70520 197350 70590
rect 197650 70520 197850 70590
rect 198150 70520 198350 70590
rect 198650 70520 198850 70590
rect 199150 70520 199350 70590
rect 199650 70520 199850 70590
rect 200150 70520 200350 70590
rect 200650 70520 200850 70590
rect 201150 70520 201350 70590
rect 201650 70520 201850 70590
rect 202150 70520 202350 70590
rect 202650 70520 202850 70590
rect 203150 70520 203350 70590
rect 203650 70520 203850 70590
rect 204150 70520 204350 70590
rect 204650 70520 204850 70590
rect 205150 70520 205350 70590
rect 205650 70520 205850 70590
rect 206150 70520 206350 70590
rect 206650 70520 206850 70590
rect 207150 70520 207350 70590
rect 207650 70520 207850 70590
rect 196150 70410 196350 70480
rect 196650 70410 196850 70480
rect 197150 70410 197350 70480
rect 197650 70410 197850 70480
rect 198150 70410 198350 70480
rect 198650 70410 198850 70480
rect 199150 70410 199350 70480
rect 199650 70410 199850 70480
rect 200150 70410 200350 70480
rect 200650 70410 200850 70480
rect 201150 70410 201350 70480
rect 201650 70410 201850 70480
rect 202150 70410 202350 70480
rect 202650 70410 202850 70480
rect 203150 70410 203350 70480
rect 203650 70410 203850 70480
rect 204150 70410 204350 70480
rect 204650 70410 204850 70480
rect 205150 70410 205350 70480
rect 205650 70410 205850 70480
rect 206150 70410 206350 70480
rect 206650 70410 206850 70480
rect 207150 70410 207350 70480
rect 207650 70410 207850 70480
rect 196020 70150 196090 70350
rect 196410 70150 196480 70350
rect 196520 70150 196590 70350
rect 196910 70150 196980 70350
rect 197020 70150 197090 70350
rect 197410 70150 197480 70350
rect 197520 70150 197590 70350
rect 197910 70150 197980 70350
rect 198020 70150 198090 70350
rect 198410 70150 198480 70350
rect 198520 70150 198590 70350
rect 198910 70150 198980 70350
rect 199020 70150 199090 70350
rect 199410 70150 199480 70350
rect 199520 70150 199590 70350
rect 199910 70150 199980 70350
rect 200020 70150 200090 70350
rect 200410 70150 200480 70350
rect 200520 70150 200590 70350
rect 200910 70150 200980 70350
rect 201020 70150 201090 70350
rect 201410 70150 201480 70350
rect 201520 70150 201590 70350
rect 201910 70150 201980 70350
rect 202020 70150 202090 70350
rect 202410 70150 202480 70350
rect 202520 70150 202590 70350
rect 202910 70150 202980 70350
rect 203020 70150 203090 70350
rect 203410 70150 203480 70350
rect 203520 70150 203590 70350
rect 203910 70150 203980 70350
rect 204020 70150 204090 70350
rect 204410 70150 204480 70350
rect 204520 70150 204590 70350
rect 204910 70150 204980 70350
rect 205020 70150 205090 70350
rect 205410 70150 205480 70350
rect 205520 70150 205590 70350
rect 205910 70150 205980 70350
rect 206020 70150 206090 70350
rect 206410 70150 206480 70350
rect 206520 70150 206590 70350
rect 206910 70150 206980 70350
rect 207020 70150 207090 70350
rect 207410 70150 207480 70350
rect 207520 70150 207590 70350
rect 207910 70150 207980 70350
rect 196150 70020 196350 70090
rect 196650 70020 196850 70090
rect 197150 70020 197350 70090
rect 197650 70020 197850 70090
rect 198150 70020 198350 70090
rect 198650 70020 198850 70090
rect 199150 70020 199350 70090
rect 199650 70020 199850 70090
rect 200150 70020 200350 70090
rect 200650 70020 200850 70090
rect 201150 70020 201350 70090
rect 201650 70020 201850 70090
rect 202150 70020 202350 70090
rect 202650 70020 202850 70090
rect 203150 70020 203350 70090
rect 203650 70020 203850 70090
rect 204150 70020 204350 70090
rect 204650 70020 204850 70090
rect 205150 70020 205350 70090
rect 205650 70020 205850 70090
rect 206150 70020 206350 70090
rect 206650 70020 206850 70090
rect 207150 70020 207350 70090
rect 207650 70020 207850 70090
rect 196150 69910 196350 69980
rect 196650 69910 196850 69980
rect 197150 69910 197350 69980
rect 197650 69910 197850 69980
rect 198150 69910 198350 69980
rect 198650 69910 198850 69980
rect 199150 69910 199350 69980
rect 199650 69910 199850 69980
rect 200150 69910 200350 69980
rect 200650 69910 200850 69980
rect 201150 69910 201350 69980
rect 201650 69910 201850 69980
rect 202150 69910 202350 69980
rect 202650 69910 202850 69980
rect 203150 69910 203350 69980
rect 203650 69910 203850 69980
rect 204150 69910 204350 69980
rect 204650 69910 204850 69980
rect 205150 69910 205350 69980
rect 205650 69910 205850 69980
rect 206150 69910 206350 69980
rect 206650 69910 206850 69980
rect 207150 69910 207350 69980
rect 207650 69910 207850 69980
rect 196020 69650 196090 69850
rect 196410 69650 196480 69850
rect 196520 69650 196590 69850
rect 196910 69650 196980 69850
rect 197020 69650 197090 69850
rect 197410 69650 197480 69850
rect 197520 69650 197590 69850
rect 197910 69650 197980 69850
rect 198020 69650 198090 69850
rect 198410 69650 198480 69850
rect 198520 69650 198590 69850
rect 198910 69650 198980 69850
rect 199020 69650 199090 69850
rect 199410 69650 199480 69850
rect 199520 69650 199590 69850
rect 199910 69650 199980 69850
rect 200020 69650 200090 69850
rect 200410 69650 200480 69850
rect 200520 69650 200590 69850
rect 200910 69650 200980 69850
rect 201020 69650 201090 69850
rect 201410 69650 201480 69850
rect 201520 69650 201590 69850
rect 201910 69650 201980 69850
rect 202020 69650 202090 69850
rect 202410 69650 202480 69850
rect 202520 69650 202590 69850
rect 202910 69650 202980 69850
rect 203020 69650 203090 69850
rect 203410 69650 203480 69850
rect 203520 69650 203590 69850
rect 203910 69650 203980 69850
rect 204020 69650 204090 69850
rect 204410 69650 204480 69850
rect 204520 69650 204590 69850
rect 204910 69650 204980 69850
rect 205020 69650 205090 69850
rect 205410 69650 205480 69850
rect 205520 69650 205590 69850
rect 205910 69650 205980 69850
rect 206020 69650 206090 69850
rect 206410 69650 206480 69850
rect 206520 69650 206590 69850
rect 206910 69650 206980 69850
rect 207020 69650 207090 69850
rect 207410 69650 207480 69850
rect 207520 69650 207590 69850
rect 207910 69650 207980 69850
rect 196150 69520 196350 69590
rect 196650 69520 196850 69590
rect 197150 69520 197350 69590
rect 197650 69520 197850 69590
rect 198150 69520 198350 69590
rect 198650 69520 198850 69590
rect 199150 69520 199350 69590
rect 199650 69520 199850 69590
rect 200150 69520 200350 69590
rect 200650 69520 200850 69590
rect 201150 69520 201350 69590
rect 201650 69520 201850 69590
rect 202150 69520 202350 69590
rect 202650 69520 202850 69590
rect 203150 69520 203350 69590
rect 203650 69520 203850 69590
rect 204150 69520 204350 69590
rect 204650 69520 204850 69590
rect 205150 69520 205350 69590
rect 205650 69520 205850 69590
rect 206150 69520 206350 69590
rect 206650 69520 206850 69590
rect 207150 69520 207350 69590
rect 207650 69520 207850 69590
rect 196150 69410 196350 69480
rect 196650 69410 196850 69480
rect 197150 69410 197350 69480
rect 197650 69410 197850 69480
rect 198150 69410 198350 69480
rect 198650 69410 198850 69480
rect 199150 69410 199350 69480
rect 199650 69410 199850 69480
rect 200150 69410 200350 69480
rect 200650 69410 200850 69480
rect 201150 69410 201350 69480
rect 201650 69410 201850 69480
rect 202150 69410 202350 69480
rect 202650 69410 202850 69480
rect 203150 69410 203350 69480
rect 203650 69410 203850 69480
rect 204150 69410 204350 69480
rect 204650 69410 204850 69480
rect 205150 69410 205350 69480
rect 205650 69410 205850 69480
rect 206150 69410 206350 69480
rect 206650 69410 206850 69480
rect 207150 69410 207350 69480
rect 207650 69410 207850 69480
rect 196020 69150 196090 69350
rect 196410 69150 196480 69350
rect 196520 69150 196590 69350
rect 196910 69150 196980 69350
rect 197020 69150 197090 69350
rect 197410 69150 197480 69350
rect 197520 69150 197590 69350
rect 197910 69150 197980 69350
rect 198020 69150 198090 69350
rect 198410 69150 198480 69350
rect 198520 69150 198590 69350
rect 198910 69150 198980 69350
rect 199020 69150 199090 69350
rect 199410 69150 199480 69350
rect 199520 69150 199590 69350
rect 199910 69150 199980 69350
rect 200020 69150 200090 69350
rect 200410 69150 200480 69350
rect 200520 69150 200590 69350
rect 200910 69150 200980 69350
rect 201020 69150 201090 69350
rect 201410 69150 201480 69350
rect 201520 69150 201590 69350
rect 201910 69150 201980 69350
rect 202020 69150 202090 69350
rect 202410 69150 202480 69350
rect 202520 69150 202590 69350
rect 202910 69150 202980 69350
rect 203020 69150 203090 69350
rect 203410 69150 203480 69350
rect 203520 69150 203590 69350
rect 203910 69150 203980 69350
rect 204020 69150 204090 69350
rect 204410 69150 204480 69350
rect 204520 69150 204590 69350
rect 204910 69150 204980 69350
rect 205020 69150 205090 69350
rect 205410 69150 205480 69350
rect 205520 69150 205590 69350
rect 205910 69150 205980 69350
rect 206020 69150 206090 69350
rect 206410 69150 206480 69350
rect 206520 69150 206590 69350
rect 206910 69150 206980 69350
rect 207020 69150 207090 69350
rect 207410 69150 207480 69350
rect 207520 69150 207590 69350
rect 207910 69150 207980 69350
rect 196150 69020 196350 69090
rect 196650 69020 196850 69090
rect 197150 69020 197350 69090
rect 197650 69020 197850 69090
rect 198150 69020 198350 69090
rect 198650 69020 198850 69090
rect 199150 69020 199350 69090
rect 199650 69020 199850 69090
rect 200150 69020 200350 69090
rect 200650 69020 200850 69090
rect 201150 69020 201350 69090
rect 201650 69020 201850 69090
rect 202150 69020 202350 69090
rect 202650 69020 202850 69090
rect 203150 69020 203350 69090
rect 203650 69020 203850 69090
rect 204150 69020 204350 69090
rect 204650 69020 204850 69090
rect 205150 69020 205350 69090
rect 205650 69020 205850 69090
rect 206150 69020 206350 69090
rect 206650 69020 206850 69090
rect 207150 69020 207350 69090
rect 207650 69020 207850 69090
rect 196150 68910 196350 68980
rect 196650 68910 196850 68980
rect 197150 68910 197350 68980
rect 197650 68910 197850 68980
rect 198150 68910 198350 68980
rect 198650 68910 198850 68980
rect 199150 68910 199350 68980
rect 199650 68910 199850 68980
rect 200150 68910 200350 68980
rect 200650 68910 200850 68980
rect 201150 68910 201350 68980
rect 201650 68910 201850 68980
rect 202150 68910 202350 68980
rect 202650 68910 202850 68980
rect 203150 68910 203350 68980
rect 203650 68910 203850 68980
rect 204150 68910 204350 68980
rect 204650 68910 204850 68980
rect 205150 68910 205350 68980
rect 205650 68910 205850 68980
rect 206150 68910 206350 68980
rect 206650 68910 206850 68980
rect 207150 68910 207350 68980
rect 207650 68910 207850 68980
rect 196020 68650 196090 68850
rect 196410 68650 196480 68850
rect 196520 68650 196590 68850
rect 196910 68650 196980 68850
rect 197020 68650 197090 68850
rect 197410 68650 197480 68850
rect 197520 68650 197590 68850
rect 197910 68650 197980 68850
rect 198020 68650 198090 68850
rect 198410 68650 198480 68850
rect 198520 68650 198590 68850
rect 198910 68650 198980 68850
rect 199020 68650 199090 68850
rect 199410 68650 199480 68850
rect 199520 68650 199590 68850
rect 199910 68650 199980 68850
rect 200020 68650 200090 68850
rect 200410 68650 200480 68850
rect 200520 68650 200590 68850
rect 200910 68650 200980 68850
rect 201020 68650 201090 68850
rect 201410 68650 201480 68850
rect 201520 68650 201590 68850
rect 201910 68650 201980 68850
rect 202020 68650 202090 68850
rect 202410 68650 202480 68850
rect 202520 68650 202590 68850
rect 202910 68650 202980 68850
rect 203020 68650 203090 68850
rect 203410 68650 203480 68850
rect 203520 68650 203590 68850
rect 203910 68650 203980 68850
rect 204020 68650 204090 68850
rect 204410 68650 204480 68850
rect 204520 68650 204590 68850
rect 204910 68650 204980 68850
rect 205020 68650 205090 68850
rect 205410 68650 205480 68850
rect 205520 68650 205590 68850
rect 205910 68650 205980 68850
rect 206020 68650 206090 68850
rect 206410 68650 206480 68850
rect 206520 68650 206590 68850
rect 206910 68650 206980 68850
rect 207020 68650 207090 68850
rect 207410 68650 207480 68850
rect 207520 68650 207590 68850
rect 207910 68650 207980 68850
rect 196150 68520 196350 68590
rect 196650 68520 196850 68590
rect 197150 68520 197350 68590
rect 197650 68520 197850 68590
rect 198150 68520 198350 68590
rect 198650 68520 198850 68590
rect 199150 68520 199350 68590
rect 199650 68520 199850 68590
rect 200150 68520 200350 68590
rect 200650 68520 200850 68590
rect 201150 68520 201350 68590
rect 201650 68520 201850 68590
rect 202150 68520 202350 68590
rect 202650 68520 202850 68590
rect 203150 68520 203350 68590
rect 203650 68520 203850 68590
rect 204150 68520 204350 68590
rect 204650 68520 204850 68590
rect 205150 68520 205350 68590
rect 205650 68520 205850 68590
rect 206150 68520 206350 68590
rect 206650 68520 206850 68590
rect 207150 68520 207350 68590
rect 207650 68520 207850 68590
rect 196150 68410 196350 68480
rect 196650 68410 196850 68480
rect 197150 68410 197350 68480
rect 197650 68410 197850 68480
rect 198150 68410 198350 68480
rect 198650 68410 198850 68480
rect 199150 68410 199350 68480
rect 199650 68410 199850 68480
rect 200150 68410 200350 68480
rect 200650 68410 200850 68480
rect 201150 68410 201350 68480
rect 201650 68410 201850 68480
rect 202150 68410 202350 68480
rect 202650 68410 202850 68480
rect 203150 68410 203350 68480
rect 203650 68410 203850 68480
rect 204150 68410 204350 68480
rect 204650 68410 204850 68480
rect 205150 68410 205350 68480
rect 205650 68410 205850 68480
rect 206150 68410 206350 68480
rect 206650 68410 206850 68480
rect 207150 68410 207350 68480
rect 207650 68410 207850 68480
rect 196020 68150 196090 68350
rect 196410 68150 196480 68350
rect 196520 68150 196590 68350
rect 196910 68150 196980 68350
rect 197020 68150 197090 68350
rect 197410 68150 197480 68350
rect 197520 68150 197590 68350
rect 197910 68150 197980 68350
rect 198020 68150 198090 68350
rect 198410 68150 198480 68350
rect 198520 68150 198590 68350
rect 198910 68150 198980 68350
rect 199020 68150 199090 68350
rect 199410 68150 199480 68350
rect 199520 68150 199590 68350
rect 199910 68150 199980 68350
rect 200020 68150 200090 68350
rect 200410 68150 200480 68350
rect 200520 68150 200590 68350
rect 200910 68150 200980 68350
rect 201020 68150 201090 68350
rect 201410 68150 201480 68350
rect 201520 68150 201590 68350
rect 201910 68150 201980 68350
rect 202020 68150 202090 68350
rect 202410 68150 202480 68350
rect 202520 68150 202590 68350
rect 202910 68150 202980 68350
rect 203020 68150 203090 68350
rect 203410 68150 203480 68350
rect 203520 68150 203590 68350
rect 203910 68150 203980 68350
rect 204020 68150 204090 68350
rect 204410 68150 204480 68350
rect 204520 68150 204590 68350
rect 204910 68150 204980 68350
rect 205020 68150 205090 68350
rect 205410 68150 205480 68350
rect 205520 68150 205590 68350
rect 205910 68150 205980 68350
rect 206020 68150 206090 68350
rect 206410 68150 206480 68350
rect 206520 68150 206590 68350
rect 206910 68150 206980 68350
rect 207020 68150 207090 68350
rect 207410 68150 207480 68350
rect 207520 68150 207590 68350
rect 207910 68150 207980 68350
rect 196150 68020 196350 68090
rect 196650 68020 196850 68090
rect 197150 68020 197350 68090
rect 197650 68020 197850 68090
rect 198150 68020 198350 68090
rect 198650 68020 198850 68090
rect 199150 68020 199350 68090
rect 199650 68020 199850 68090
rect 200150 68020 200350 68090
rect 200650 68020 200850 68090
rect 201150 68020 201350 68090
rect 201650 68020 201850 68090
rect 202150 68020 202350 68090
rect 202650 68020 202850 68090
rect 203150 68020 203350 68090
rect 203650 68020 203850 68090
rect 204150 68020 204350 68090
rect 204650 68020 204850 68090
rect 205150 68020 205350 68090
rect 205650 68020 205850 68090
rect 206150 68020 206350 68090
rect 206650 68020 206850 68090
rect 207150 68020 207350 68090
rect 207650 68020 207850 68090
rect 196150 67910 196350 67980
rect 196650 67910 196850 67980
rect 197150 67910 197350 67980
rect 197650 67910 197850 67980
rect 198150 67910 198350 67980
rect 198650 67910 198850 67980
rect 199150 67910 199350 67980
rect 199650 67910 199850 67980
rect 200150 67910 200350 67980
rect 200650 67910 200850 67980
rect 201150 67910 201350 67980
rect 201650 67910 201850 67980
rect 202150 67910 202350 67980
rect 202650 67910 202850 67980
rect 203150 67910 203350 67980
rect 203650 67910 203850 67980
rect 204150 67910 204350 67980
rect 204650 67910 204850 67980
rect 205150 67910 205350 67980
rect 205650 67910 205850 67980
rect 206150 67910 206350 67980
rect 206650 67910 206850 67980
rect 207150 67910 207350 67980
rect 207650 67910 207850 67980
rect 196020 67650 196090 67850
rect 196410 67650 196480 67850
rect 196520 67650 196590 67850
rect 196910 67650 196980 67850
rect 197020 67650 197090 67850
rect 197410 67650 197480 67850
rect 197520 67650 197590 67850
rect 197910 67650 197980 67850
rect 198020 67650 198090 67850
rect 198410 67650 198480 67850
rect 198520 67650 198590 67850
rect 198910 67650 198980 67850
rect 199020 67650 199090 67850
rect 199410 67650 199480 67850
rect 199520 67650 199590 67850
rect 199910 67650 199980 67850
rect 200020 67650 200090 67850
rect 200410 67650 200480 67850
rect 200520 67650 200590 67850
rect 200910 67650 200980 67850
rect 201020 67650 201090 67850
rect 201410 67650 201480 67850
rect 201520 67650 201590 67850
rect 201910 67650 201980 67850
rect 202020 67650 202090 67850
rect 202410 67650 202480 67850
rect 202520 67650 202590 67850
rect 202910 67650 202980 67850
rect 203020 67650 203090 67850
rect 203410 67650 203480 67850
rect 203520 67650 203590 67850
rect 203910 67650 203980 67850
rect 204020 67650 204090 67850
rect 204410 67650 204480 67850
rect 204520 67650 204590 67850
rect 204910 67650 204980 67850
rect 205020 67650 205090 67850
rect 205410 67650 205480 67850
rect 205520 67650 205590 67850
rect 205910 67650 205980 67850
rect 206020 67650 206090 67850
rect 206410 67650 206480 67850
rect 206520 67650 206590 67850
rect 206910 67650 206980 67850
rect 207020 67650 207090 67850
rect 207410 67650 207480 67850
rect 207520 67650 207590 67850
rect 207910 67650 207980 67850
rect 196150 67520 196350 67590
rect 196650 67520 196850 67590
rect 197150 67520 197350 67590
rect 197650 67520 197850 67590
rect 198150 67520 198350 67590
rect 198650 67520 198850 67590
rect 199150 67520 199350 67590
rect 199650 67520 199850 67590
rect 200150 67520 200350 67590
rect 200650 67520 200850 67590
rect 201150 67520 201350 67590
rect 201650 67520 201850 67590
rect 202150 67520 202350 67590
rect 202650 67520 202850 67590
rect 203150 67520 203350 67590
rect 203650 67520 203850 67590
rect 204150 67520 204350 67590
rect 204650 67520 204850 67590
rect 205150 67520 205350 67590
rect 205650 67520 205850 67590
rect 206150 67520 206350 67590
rect 206650 67520 206850 67590
rect 207150 67520 207350 67590
rect 207650 67520 207850 67590
rect 196150 67410 196350 67480
rect 196650 67410 196850 67480
rect 197150 67410 197350 67480
rect 197650 67410 197850 67480
rect 198150 67410 198350 67480
rect 198650 67410 198850 67480
rect 199150 67410 199350 67480
rect 199650 67410 199850 67480
rect 200150 67410 200350 67480
rect 200650 67410 200850 67480
rect 201150 67410 201350 67480
rect 201650 67410 201850 67480
rect 202150 67410 202350 67480
rect 202650 67410 202850 67480
rect 203150 67410 203350 67480
rect 203650 67410 203850 67480
rect 204150 67410 204350 67480
rect 204650 67410 204850 67480
rect 205150 67410 205350 67480
rect 205650 67410 205850 67480
rect 206150 67410 206350 67480
rect 206650 67410 206850 67480
rect 207150 67410 207350 67480
rect 207650 67410 207850 67480
rect 196020 67150 196090 67350
rect 196410 67150 196480 67350
rect 196520 67150 196590 67350
rect 196910 67150 196980 67350
rect 197020 67150 197090 67350
rect 197410 67150 197480 67350
rect 197520 67150 197590 67350
rect 197910 67150 197980 67350
rect 198020 67150 198090 67350
rect 198410 67150 198480 67350
rect 198520 67150 198590 67350
rect 198910 67150 198980 67350
rect 199020 67150 199090 67350
rect 199410 67150 199480 67350
rect 199520 67150 199590 67350
rect 199910 67150 199980 67350
rect 200020 67150 200090 67350
rect 200410 67150 200480 67350
rect 200520 67150 200590 67350
rect 200910 67150 200980 67350
rect 201020 67150 201090 67350
rect 201410 67150 201480 67350
rect 201520 67150 201590 67350
rect 201910 67150 201980 67350
rect 202020 67150 202090 67350
rect 202410 67150 202480 67350
rect 202520 67150 202590 67350
rect 202910 67150 202980 67350
rect 203020 67150 203090 67350
rect 203410 67150 203480 67350
rect 203520 67150 203590 67350
rect 203910 67150 203980 67350
rect 204020 67150 204090 67350
rect 204410 67150 204480 67350
rect 204520 67150 204590 67350
rect 204910 67150 204980 67350
rect 205020 67150 205090 67350
rect 205410 67150 205480 67350
rect 205520 67150 205590 67350
rect 205910 67150 205980 67350
rect 206020 67150 206090 67350
rect 206410 67150 206480 67350
rect 206520 67150 206590 67350
rect 206910 67150 206980 67350
rect 207020 67150 207090 67350
rect 207410 67150 207480 67350
rect 207520 67150 207590 67350
rect 207910 67150 207980 67350
rect 196150 67020 196350 67090
rect 196650 67020 196850 67090
rect 197150 67020 197350 67090
rect 197650 67020 197850 67090
rect 198150 67020 198350 67090
rect 198650 67020 198850 67090
rect 199150 67020 199350 67090
rect 199650 67020 199850 67090
rect 200150 67020 200350 67090
rect 200650 67020 200850 67090
rect 201150 67020 201350 67090
rect 201650 67020 201850 67090
rect 202150 67020 202350 67090
rect 202650 67020 202850 67090
rect 203150 67020 203350 67090
rect 203650 67020 203850 67090
rect 204150 67020 204350 67090
rect 204650 67020 204850 67090
rect 205150 67020 205350 67090
rect 205650 67020 205850 67090
rect 206150 67020 206350 67090
rect 206650 67020 206850 67090
rect 207150 67020 207350 67090
rect 207650 67020 207850 67090
rect 196150 66910 196350 66980
rect 196650 66910 196850 66980
rect 197150 66910 197350 66980
rect 197650 66910 197850 66980
rect 198150 66910 198350 66980
rect 198650 66910 198850 66980
rect 199150 66910 199350 66980
rect 199650 66910 199850 66980
rect 200150 66910 200350 66980
rect 200650 66910 200850 66980
rect 201150 66910 201350 66980
rect 201650 66910 201850 66980
rect 202150 66910 202350 66980
rect 202650 66910 202850 66980
rect 203150 66910 203350 66980
rect 203650 66910 203850 66980
rect 204150 66910 204350 66980
rect 204650 66910 204850 66980
rect 205150 66910 205350 66980
rect 205650 66910 205850 66980
rect 206150 66910 206350 66980
rect 206650 66910 206850 66980
rect 207150 66910 207350 66980
rect 207650 66910 207850 66980
rect 196020 66650 196090 66850
rect 196410 66650 196480 66850
rect 196520 66650 196590 66850
rect 196910 66650 196980 66850
rect 197020 66650 197090 66850
rect 197410 66650 197480 66850
rect 197520 66650 197590 66850
rect 197910 66650 197980 66850
rect 198020 66650 198090 66850
rect 198410 66650 198480 66850
rect 198520 66650 198590 66850
rect 198910 66650 198980 66850
rect 199020 66650 199090 66850
rect 199410 66650 199480 66850
rect 199520 66650 199590 66850
rect 199910 66650 199980 66850
rect 200020 66650 200090 66850
rect 200410 66650 200480 66850
rect 200520 66650 200590 66850
rect 200910 66650 200980 66850
rect 201020 66650 201090 66850
rect 201410 66650 201480 66850
rect 201520 66650 201590 66850
rect 201910 66650 201980 66850
rect 202020 66650 202090 66850
rect 202410 66650 202480 66850
rect 202520 66650 202590 66850
rect 202910 66650 202980 66850
rect 203020 66650 203090 66850
rect 203410 66650 203480 66850
rect 203520 66650 203590 66850
rect 203910 66650 203980 66850
rect 204020 66650 204090 66850
rect 204410 66650 204480 66850
rect 204520 66650 204590 66850
rect 204910 66650 204980 66850
rect 205020 66650 205090 66850
rect 205410 66650 205480 66850
rect 205520 66650 205590 66850
rect 205910 66650 205980 66850
rect 206020 66650 206090 66850
rect 206410 66650 206480 66850
rect 206520 66650 206590 66850
rect 206910 66650 206980 66850
rect 207020 66650 207090 66850
rect 207410 66650 207480 66850
rect 207520 66650 207590 66850
rect 207910 66650 207980 66850
rect 196150 66520 196350 66590
rect 196650 66520 196850 66590
rect 197150 66520 197350 66590
rect 197650 66520 197850 66590
rect 198150 66520 198350 66590
rect 198650 66520 198850 66590
rect 199150 66520 199350 66590
rect 199650 66520 199850 66590
rect 200150 66520 200350 66590
rect 200650 66520 200850 66590
rect 201150 66520 201350 66590
rect 201650 66520 201850 66590
rect 202150 66520 202350 66590
rect 202650 66520 202850 66590
rect 203150 66520 203350 66590
rect 203650 66520 203850 66590
rect 204150 66520 204350 66590
rect 204650 66520 204850 66590
rect 205150 66520 205350 66590
rect 205650 66520 205850 66590
rect 206150 66520 206350 66590
rect 206650 66520 206850 66590
rect 207150 66520 207350 66590
rect 207650 66520 207850 66590
rect 196150 66410 196350 66480
rect 196650 66410 196850 66480
rect 197150 66410 197350 66480
rect 197650 66410 197850 66480
rect 198150 66410 198350 66480
rect 198650 66410 198850 66480
rect 199150 66410 199350 66480
rect 199650 66410 199850 66480
rect 200150 66410 200350 66480
rect 200650 66410 200850 66480
rect 201150 66410 201350 66480
rect 201650 66410 201850 66480
rect 202150 66410 202350 66480
rect 202650 66410 202850 66480
rect 203150 66410 203350 66480
rect 203650 66410 203850 66480
rect 204150 66410 204350 66480
rect 204650 66410 204850 66480
rect 205150 66410 205350 66480
rect 205650 66410 205850 66480
rect 206150 66410 206350 66480
rect 206650 66410 206850 66480
rect 207150 66410 207350 66480
rect 207650 66410 207850 66480
rect 196020 66150 196090 66350
rect 196410 66150 196480 66350
rect 196520 66150 196590 66350
rect 196910 66150 196980 66350
rect 197020 66150 197090 66350
rect 197410 66150 197480 66350
rect 197520 66150 197590 66350
rect 197910 66150 197980 66350
rect 198020 66150 198090 66350
rect 198410 66150 198480 66350
rect 198520 66150 198590 66350
rect 198910 66150 198980 66350
rect 199020 66150 199090 66350
rect 199410 66150 199480 66350
rect 199520 66150 199590 66350
rect 199910 66150 199980 66350
rect 200020 66150 200090 66350
rect 200410 66150 200480 66350
rect 200520 66150 200590 66350
rect 200910 66150 200980 66350
rect 201020 66150 201090 66350
rect 201410 66150 201480 66350
rect 201520 66150 201590 66350
rect 201910 66150 201980 66350
rect 202020 66150 202090 66350
rect 202410 66150 202480 66350
rect 202520 66150 202590 66350
rect 202910 66150 202980 66350
rect 203020 66150 203090 66350
rect 203410 66150 203480 66350
rect 203520 66150 203590 66350
rect 203910 66150 203980 66350
rect 204020 66150 204090 66350
rect 204410 66150 204480 66350
rect 204520 66150 204590 66350
rect 204910 66150 204980 66350
rect 205020 66150 205090 66350
rect 205410 66150 205480 66350
rect 205520 66150 205590 66350
rect 205910 66150 205980 66350
rect 206020 66150 206090 66350
rect 206410 66150 206480 66350
rect 206520 66150 206590 66350
rect 206910 66150 206980 66350
rect 207020 66150 207090 66350
rect 207410 66150 207480 66350
rect 207520 66150 207590 66350
rect 207910 66150 207980 66350
rect 196150 66020 196350 66090
rect 196650 66020 196850 66090
rect 197150 66020 197350 66090
rect 197650 66020 197850 66090
rect 198150 66020 198350 66090
rect 198650 66020 198850 66090
rect 199150 66020 199350 66090
rect 199650 66020 199850 66090
rect 200150 66020 200350 66090
rect 200650 66020 200850 66090
rect 201150 66020 201350 66090
rect 201650 66020 201850 66090
rect 202150 66020 202350 66090
rect 202650 66020 202850 66090
rect 203150 66020 203350 66090
rect 203650 66020 203850 66090
rect 204150 66020 204350 66090
rect 204650 66020 204850 66090
rect 205150 66020 205350 66090
rect 205650 66020 205850 66090
rect 206150 66020 206350 66090
rect 206650 66020 206850 66090
rect 207150 66020 207350 66090
rect 207650 66020 207850 66090
rect 190150 65910 190350 65980
rect 190650 65910 190850 65980
rect 191150 65910 191350 65980
rect 191650 65910 191850 65980
rect 192150 65910 192350 65980
rect 192650 65910 192850 65980
rect 193150 65910 193350 65980
rect 193650 65910 193850 65980
rect 194150 65910 194350 65980
rect 194650 65910 194850 65980
rect 195150 65910 195350 65980
rect 195650 65910 195850 65980
rect 196150 65910 196350 65980
rect 196650 65910 196850 65980
rect 197150 65910 197350 65980
rect 197650 65910 197850 65980
rect 198150 65910 198350 65980
rect 198650 65910 198850 65980
rect 199150 65910 199350 65980
rect 199650 65910 199850 65980
rect 200150 65910 200350 65980
rect 200650 65910 200850 65980
rect 201150 65910 201350 65980
rect 201650 65910 201850 65980
rect 202150 65910 202350 65980
rect 202650 65910 202850 65980
rect 203150 65910 203350 65980
rect 203650 65910 203850 65980
rect 204150 65910 204350 65980
rect 204650 65910 204850 65980
rect 205150 65910 205350 65980
rect 205650 65910 205850 65980
rect 206150 65910 206350 65980
rect 206650 65910 206850 65980
rect 207150 65910 207350 65980
rect 207650 65910 207850 65980
rect 190020 65650 190090 65850
rect 190410 65650 190480 65850
rect 190520 65650 190590 65850
rect 190910 65650 190980 65850
rect 191020 65650 191090 65850
rect 191410 65650 191480 65850
rect 191520 65650 191590 65850
rect 191910 65650 191980 65850
rect 192020 65650 192090 65850
rect 192410 65650 192480 65850
rect 192520 65650 192590 65850
rect 192910 65650 192980 65850
rect 193020 65650 193090 65850
rect 193410 65650 193480 65850
rect 193520 65650 193590 65850
rect 193910 65650 193980 65850
rect 194020 65650 194090 65850
rect 194410 65650 194480 65850
rect 194520 65650 194590 65850
rect 194910 65650 194980 65850
rect 195020 65650 195090 65850
rect 195410 65650 195480 65850
rect 195520 65650 195590 65850
rect 195910 65650 195980 65850
rect 196020 65650 196090 65850
rect 196410 65650 196480 65850
rect 196520 65650 196590 65850
rect 196910 65650 196980 65850
rect 197020 65650 197090 65850
rect 197410 65650 197480 65850
rect 197520 65650 197590 65850
rect 197910 65650 197980 65850
rect 198020 65650 198090 65850
rect 198410 65650 198480 65850
rect 198520 65650 198590 65850
rect 198910 65650 198980 65850
rect 199020 65650 199090 65850
rect 199410 65650 199480 65850
rect 199520 65650 199590 65850
rect 199910 65650 199980 65850
rect 200020 65650 200090 65850
rect 200410 65650 200480 65850
rect 200520 65650 200590 65850
rect 200910 65650 200980 65850
rect 201020 65650 201090 65850
rect 201410 65650 201480 65850
rect 201520 65650 201590 65850
rect 201910 65650 201980 65850
rect 202020 65650 202090 65850
rect 202410 65650 202480 65850
rect 202520 65650 202590 65850
rect 202910 65650 202980 65850
rect 203020 65650 203090 65850
rect 203410 65650 203480 65850
rect 203520 65650 203590 65850
rect 203910 65650 203980 65850
rect 204020 65650 204090 65850
rect 204410 65650 204480 65850
rect 204520 65650 204590 65850
rect 204910 65650 204980 65850
rect 205020 65650 205090 65850
rect 205410 65650 205480 65850
rect 205520 65650 205590 65850
rect 205910 65650 205980 65850
rect 206020 65650 206090 65850
rect 206410 65650 206480 65850
rect 206520 65650 206590 65850
rect 206910 65650 206980 65850
rect 207020 65650 207090 65850
rect 207410 65650 207480 65850
rect 207520 65650 207590 65850
rect 207910 65650 207980 65850
rect 190150 65520 190350 65590
rect 190650 65520 190850 65590
rect 191150 65520 191350 65590
rect 191650 65520 191850 65590
rect 192150 65520 192350 65590
rect 192650 65520 192850 65590
rect 193150 65520 193350 65590
rect 193650 65520 193850 65590
rect 194150 65520 194350 65590
rect 194650 65520 194850 65590
rect 195150 65520 195350 65590
rect 195650 65520 195850 65590
rect 196150 65520 196350 65590
rect 196650 65520 196850 65590
rect 197150 65520 197350 65590
rect 197650 65520 197850 65590
rect 198150 65520 198350 65590
rect 198650 65520 198850 65590
rect 199150 65520 199350 65590
rect 199650 65520 199850 65590
rect 200150 65520 200350 65590
rect 200650 65520 200850 65590
rect 201150 65520 201350 65590
rect 201650 65520 201850 65590
rect 202150 65520 202350 65590
rect 202650 65520 202850 65590
rect 203150 65520 203350 65590
rect 203650 65520 203850 65590
rect 204150 65520 204350 65590
rect 204650 65520 204850 65590
rect 205150 65520 205350 65590
rect 205650 65520 205850 65590
rect 206150 65520 206350 65590
rect 206650 65520 206850 65590
rect 207150 65520 207350 65590
rect 207650 65520 207850 65590
rect 190150 65410 190350 65480
rect 190650 65410 190850 65480
rect 191150 65410 191350 65480
rect 191650 65410 191850 65480
rect 192150 65410 192350 65480
rect 192650 65410 192850 65480
rect 193150 65410 193350 65480
rect 193650 65410 193850 65480
rect 194150 65410 194350 65480
rect 194650 65410 194850 65480
rect 195150 65410 195350 65480
rect 195650 65410 195850 65480
rect 196150 65410 196350 65480
rect 196650 65410 196850 65480
rect 197150 65410 197350 65480
rect 197650 65410 197850 65480
rect 198150 65410 198350 65480
rect 198650 65410 198850 65480
rect 199150 65410 199350 65480
rect 199650 65410 199850 65480
rect 200150 65410 200350 65480
rect 200650 65410 200850 65480
rect 201150 65410 201350 65480
rect 201650 65410 201850 65480
rect 202150 65410 202350 65480
rect 202650 65410 202850 65480
rect 203150 65410 203350 65480
rect 203650 65410 203850 65480
rect 204150 65410 204350 65480
rect 204650 65410 204850 65480
rect 205150 65410 205350 65480
rect 205650 65410 205850 65480
rect 206150 65410 206350 65480
rect 206650 65410 206850 65480
rect 207150 65410 207350 65480
rect 207650 65410 207850 65480
rect 190020 65150 190090 65350
rect 190410 65150 190480 65350
rect 190520 65150 190590 65350
rect 190910 65150 190980 65350
rect 191020 65150 191090 65350
rect 191410 65150 191480 65350
rect 191520 65150 191590 65350
rect 191910 65150 191980 65350
rect 192020 65150 192090 65350
rect 192410 65150 192480 65350
rect 192520 65150 192590 65350
rect 192910 65150 192980 65350
rect 193020 65150 193090 65350
rect 193410 65150 193480 65350
rect 193520 65150 193590 65350
rect 193910 65150 193980 65350
rect 194020 65150 194090 65350
rect 194410 65150 194480 65350
rect 194520 65150 194590 65350
rect 194910 65150 194980 65350
rect 195020 65150 195090 65350
rect 195410 65150 195480 65350
rect 195520 65150 195590 65350
rect 195910 65150 195980 65350
rect 196020 65150 196090 65350
rect 196410 65150 196480 65350
rect 196520 65150 196590 65350
rect 196910 65150 196980 65350
rect 197020 65150 197090 65350
rect 197410 65150 197480 65350
rect 197520 65150 197590 65350
rect 197910 65150 197980 65350
rect 198020 65150 198090 65350
rect 198410 65150 198480 65350
rect 198520 65150 198590 65350
rect 198910 65150 198980 65350
rect 199020 65150 199090 65350
rect 199410 65150 199480 65350
rect 199520 65150 199590 65350
rect 199910 65150 199980 65350
rect 200020 65150 200090 65350
rect 200410 65150 200480 65350
rect 200520 65150 200590 65350
rect 200910 65150 200980 65350
rect 201020 65150 201090 65350
rect 201410 65150 201480 65350
rect 201520 65150 201590 65350
rect 201910 65150 201980 65350
rect 202020 65150 202090 65350
rect 202410 65150 202480 65350
rect 202520 65150 202590 65350
rect 202910 65150 202980 65350
rect 203020 65150 203090 65350
rect 203410 65150 203480 65350
rect 203520 65150 203590 65350
rect 203910 65150 203980 65350
rect 204020 65150 204090 65350
rect 204410 65150 204480 65350
rect 204520 65150 204590 65350
rect 204910 65150 204980 65350
rect 205020 65150 205090 65350
rect 205410 65150 205480 65350
rect 205520 65150 205590 65350
rect 205910 65150 205980 65350
rect 206020 65150 206090 65350
rect 206410 65150 206480 65350
rect 206520 65150 206590 65350
rect 206910 65150 206980 65350
rect 207020 65150 207090 65350
rect 207410 65150 207480 65350
rect 207520 65150 207590 65350
rect 207910 65150 207980 65350
rect 190150 65020 190350 65090
rect 190650 65020 190850 65090
rect 191150 65020 191350 65090
rect 191650 65020 191850 65090
rect 192150 65020 192350 65090
rect 192650 65020 192850 65090
rect 193150 65020 193350 65090
rect 193650 65020 193850 65090
rect 194150 65020 194350 65090
rect 194650 65020 194850 65090
rect 195150 65020 195350 65090
rect 195650 65020 195850 65090
rect 196150 65020 196350 65090
rect 196650 65020 196850 65090
rect 197150 65020 197350 65090
rect 197650 65020 197850 65090
rect 198150 65020 198350 65090
rect 198650 65020 198850 65090
rect 199150 65020 199350 65090
rect 199650 65020 199850 65090
rect 200150 65020 200350 65090
rect 200650 65020 200850 65090
rect 201150 65020 201350 65090
rect 201650 65020 201850 65090
rect 202150 65020 202350 65090
rect 202650 65020 202850 65090
rect 203150 65020 203350 65090
rect 203650 65020 203850 65090
rect 204150 65020 204350 65090
rect 204650 65020 204850 65090
rect 205150 65020 205350 65090
rect 205650 65020 205850 65090
rect 206150 65020 206350 65090
rect 206650 65020 206850 65090
rect 207150 65020 207350 65090
rect 207650 65020 207850 65090
rect 190150 64910 190350 64980
rect 190650 64910 190850 64980
rect 191150 64910 191350 64980
rect 191650 64910 191850 64980
rect 192150 64910 192350 64980
rect 192650 64910 192850 64980
rect 193150 64910 193350 64980
rect 193650 64910 193850 64980
rect 194150 64910 194350 64980
rect 194650 64910 194850 64980
rect 195150 64910 195350 64980
rect 195650 64910 195850 64980
rect 196150 64910 196350 64980
rect 196650 64910 196850 64980
rect 197150 64910 197350 64980
rect 197650 64910 197850 64980
rect 198150 64910 198350 64980
rect 198650 64910 198850 64980
rect 199150 64910 199350 64980
rect 199650 64910 199850 64980
rect 200150 64910 200350 64980
rect 200650 64910 200850 64980
rect 201150 64910 201350 64980
rect 201650 64910 201850 64980
rect 202150 64910 202350 64980
rect 202650 64910 202850 64980
rect 203150 64910 203350 64980
rect 203650 64910 203850 64980
rect 204150 64910 204350 64980
rect 204650 64910 204850 64980
rect 205150 64910 205350 64980
rect 205650 64910 205850 64980
rect 206150 64910 206350 64980
rect 206650 64910 206850 64980
rect 207150 64910 207350 64980
rect 207650 64910 207850 64980
rect 190020 64650 190090 64850
rect 190410 64650 190480 64850
rect 190520 64650 190590 64850
rect 190910 64650 190980 64850
rect 191020 64650 191090 64850
rect 191410 64650 191480 64850
rect 191520 64650 191590 64850
rect 191910 64650 191980 64850
rect 192020 64650 192090 64850
rect 192410 64650 192480 64850
rect 192520 64650 192590 64850
rect 192910 64650 192980 64850
rect 193020 64650 193090 64850
rect 193410 64650 193480 64850
rect 193520 64650 193590 64850
rect 193910 64650 193980 64850
rect 194020 64650 194090 64850
rect 194410 64650 194480 64850
rect 194520 64650 194590 64850
rect 194910 64650 194980 64850
rect 195020 64650 195090 64850
rect 195410 64650 195480 64850
rect 195520 64650 195590 64850
rect 195910 64650 195980 64850
rect 196020 64650 196090 64850
rect 196410 64650 196480 64850
rect 196520 64650 196590 64850
rect 196910 64650 196980 64850
rect 197020 64650 197090 64850
rect 197410 64650 197480 64850
rect 197520 64650 197590 64850
rect 197910 64650 197980 64850
rect 198020 64650 198090 64850
rect 198410 64650 198480 64850
rect 198520 64650 198590 64850
rect 198910 64650 198980 64850
rect 199020 64650 199090 64850
rect 199410 64650 199480 64850
rect 199520 64650 199590 64850
rect 199910 64650 199980 64850
rect 200020 64650 200090 64850
rect 200410 64650 200480 64850
rect 200520 64650 200590 64850
rect 200910 64650 200980 64850
rect 201020 64650 201090 64850
rect 201410 64650 201480 64850
rect 201520 64650 201590 64850
rect 201910 64650 201980 64850
rect 202020 64650 202090 64850
rect 202410 64650 202480 64850
rect 202520 64650 202590 64850
rect 202910 64650 202980 64850
rect 203020 64650 203090 64850
rect 203410 64650 203480 64850
rect 203520 64650 203590 64850
rect 203910 64650 203980 64850
rect 204020 64650 204090 64850
rect 204410 64650 204480 64850
rect 204520 64650 204590 64850
rect 204910 64650 204980 64850
rect 205020 64650 205090 64850
rect 205410 64650 205480 64850
rect 205520 64650 205590 64850
rect 205910 64650 205980 64850
rect 206020 64650 206090 64850
rect 206410 64650 206480 64850
rect 206520 64650 206590 64850
rect 206910 64650 206980 64850
rect 207020 64650 207090 64850
rect 207410 64650 207480 64850
rect 207520 64650 207590 64850
rect 207910 64650 207980 64850
rect 190150 64520 190350 64590
rect 190650 64520 190850 64590
rect 191150 64520 191350 64590
rect 191650 64520 191850 64590
rect 192150 64520 192350 64590
rect 192650 64520 192850 64590
rect 193150 64520 193350 64590
rect 193650 64520 193850 64590
rect 194150 64520 194350 64590
rect 194650 64520 194850 64590
rect 195150 64520 195350 64590
rect 195650 64520 195850 64590
rect 196150 64520 196350 64590
rect 196650 64520 196850 64590
rect 197150 64520 197350 64590
rect 197650 64520 197850 64590
rect 198150 64520 198350 64590
rect 198650 64520 198850 64590
rect 199150 64520 199350 64590
rect 199650 64520 199850 64590
rect 200150 64520 200350 64590
rect 200650 64520 200850 64590
rect 201150 64520 201350 64590
rect 201650 64520 201850 64590
rect 202150 64520 202350 64590
rect 202650 64520 202850 64590
rect 203150 64520 203350 64590
rect 203650 64520 203850 64590
rect 204150 64520 204350 64590
rect 204650 64520 204850 64590
rect 205150 64520 205350 64590
rect 205650 64520 205850 64590
rect 206150 64520 206350 64590
rect 206650 64520 206850 64590
rect 207150 64520 207350 64590
rect 207650 64520 207850 64590
rect 190150 64410 190350 64480
rect 190650 64410 190850 64480
rect 191150 64410 191350 64480
rect 191650 64410 191850 64480
rect 192150 64410 192350 64480
rect 192650 64410 192850 64480
rect 193150 64410 193350 64480
rect 193650 64410 193850 64480
rect 194150 64410 194350 64480
rect 194650 64410 194850 64480
rect 195150 64410 195350 64480
rect 195650 64410 195850 64480
rect 196150 64410 196350 64480
rect 196650 64410 196850 64480
rect 197150 64410 197350 64480
rect 197650 64410 197850 64480
rect 198150 64410 198350 64480
rect 198650 64410 198850 64480
rect 199150 64410 199350 64480
rect 199650 64410 199850 64480
rect 200150 64410 200350 64480
rect 200650 64410 200850 64480
rect 201150 64410 201350 64480
rect 201650 64410 201850 64480
rect 202150 64410 202350 64480
rect 202650 64410 202850 64480
rect 203150 64410 203350 64480
rect 203650 64410 203850 64480
rect 204150 64410 204350 64480
rect 204650 64410 204850 64480
rect 205150 64410 205350 64480
rect 205650 64410 205850 64480
rect 206150 64410 206350 64480
rect 206650 64410 206850 64480
rect 207150 64410 207350 64480
rect 207650 64410 207850 64480
rect 190020 64150 190090 64350
rect 190410 64150 190480 64350
rect 190520 64150 190590 64350
rect 190910 64150 190980 64350
rect 191020 64150 191090 64350
rect 191410 64150 191480 64350
rect 191520 64150 191590 64350
rect 191910 64150 191980 64350
rect 192020 64150 192090 64350
rect 192410 64150 192480 64350
rect 192520 64150 192590 64350
rect 192910 64150 192980 64350
rect 193020 64150 193090 64350
rect 193410 64150 193480 64350
rect 193520 64150 193590 64350
rect 193910 64150 193980 64350
rect 194020 64150 194090 64350
rect 194410 64150 194480 64350
rect 194520 64150 194590 64350
rect 194910 64150 194980 64350
rect 195020 64150 195090 64350
rect 195410 64150 195480 64350
rect 195520 64150 195590 64350
rect 195910 64150 195980 64350
rect 196020 64150 196090 64350
rect 196410 64150 196480 64350
rect 196520 64150 196590 64350
rect 196910 64150 196980 64350
rect 197020 64150 197090 64350
rect 197410 64150 197480 64350
rect 197520 64150 197590 64350
rect 197910 64150 197980 64350
rect 198020 64150 198090 64350
rect 198410 64150 198480 64350
rect 198520 64150 198590 64350
rect 198910 64150 198980 64350
rect 199020 64150 199090 64350
rect 199410 64150 199480 64350
rect 199520 64150 199590 64350
rect 199910 64150 199980 64350
rect 200020 64150 200090 64350
rect 200410 64150 200480 64350
rect 200520 64150 200590 64350
rect 200910 64150 200980 64350
rect 201020 64150 201090 64350
rect 201410 64150 201480 64350
rect 201520 64150 201590 64350
rect 201910 64150 201980 64350
rect 202020 64150 202090 64350
rect 202410 64150 202480 64350
rect 202520 64150 202590 64350
rect 202910 64150 202980 64350
rect 203020 64150 203090 64350
rect 203410 64150 203480 64350
rect 203520 64150 203590 64350
rect 203910 64150 203980 64350
rect 204020 64150 204090 64350
rect 204410 64150 204480 64350
rect 204520 64150 204590 64350
rect 204910 64150 204980 64350
rect 205020 64150 205090 64350
rect 205410 64150 205480 64350
rect 205520 64150 205590 64350
rect 205910 64150 205980 64350
rect 206020 64150 206090 64350
rect 206410 64150 206480 64350
rect 206520 64150 206590 64350
rect 206910 64150 206980 64350
rect 207020 64150 207090 64350
rect 207410 64150 207480 64350
rect 207520 64150 207590 64350
rect 207910 64150 207980 64350
rect 190150 64020 190350 64090
rect 190650 64020 190850 64090
rect 191150 64020 191350 64090
rect 191650 64020 191850 64090
rect 192150 64020 192350 64090
rect 192650 64020 192850 64090
rect 193150 64020 193350 64090
rect 193650 64020 193850 64090
rect 194150 64020 194350 64090
rect 194650 64020 194850 64090
rect 195150 64020 195350 64090
rect 195650 64020 195850 64090
rect 196150 64020 196350 64090
rect 196650 64020 196850 64090
rect 197150 64020 197350 64090
rect 197650 64020 197850 64090
rect 198150 64020 198350 64090
rect 198650 64020 198850 64090
rect 199150 64020 199350 64090
rect 199650 64020 199850 64090
rect 200150 64020 200350 64090
rect 200650 64020 200850 64090
rect 201150 64020 201350 64090
rect 201650 64020 201850 64090
rect 202150 64020 202350 64090
rect 202650 64020 202850 64090
rect 203150 64020 203350 64090
rect 203650 64020 203850 64090
rect 204150 64020 204350 64090
rect 204650 64020 204850 64090
rect 205150 64020 205350 64090
rect 205650 64020 205850 64090
rect 206150 64020 206350 64090
rect 206650 64020 206850 64090
rect 207150 64020 207350 64090
rect 207650 64020 207850 64090
rect 204150 63910 204350 63980
rect 204650 63910 204850 63980
rect 205150 63910 205350 63980
rect 205650 63910 205850 63980
rect 206150 63910 206350 63980
rect 206650 63910 206850 63980
rect 207150 63910 207350 63980
rect 207650 63910 207850 63980
rect 204020 63650 204090 63850
rect 204410 63650 204480 63850
rect 204520 63650 204590 63850
rect 204910 63650 204980 63850
rect 205020 63650 205090 63850
rect 205410 63650 205480 63850
rect 205520 63650 205590 63850
rect 205910 63650 205980 63850
rect 206020 63650 206090 63850
rect 206410 63650 206480 63850
rect 206520 63650 206590 63850
rect 206910 63650 206980 63850
rect 207020 63650 207090 63850
rect 207410 63650 207480 63850
rect 207520 63650 207590 63850
rect 207910 63650 207980 63850
rect 204150 63520 204350 63590
rect 204650 63520 204850 63590
rect 205150 63520 205350 63590
rect 205650 63520 205850 63590
rect 206150 63520 206350 63590
rect 206650 63520 206850 63590
rect 207150 63520 207350 63590
rect 207650 63520 207850 63590
rect 204150 63410 204350 63480
rect 204650 63410 204850 63480
rect 205150 63410 205350 63480
rect 205650 63410 205850 63480
rect 206150 63410 206350 63480
rect 206650 63410 206850 63480
rect 207150 63410 207350 63480
rect 207650 63410 207850 63480
rect 204020 63150 204090 63350
rect 204410 63150 204480 63350
rect 204520 63150 204590 63350
rect 204910 63150 204980 63350
rect 205020 63150 205090 63350
rect 205410 63150 205480 63350
rect 205520 63150 205590 63350
rect 205910 63150 205980 63350
rect 206020 63150 206090 63350
rect 206410 63150 206480 63350
rect 206520 63150 206590 63350
rect 206910 63150 206980 63350
rect 207020 63150 207090 63350
rect 207410 63150 207480 63350
rect 207520 63150 207590 63350
rect 207910 63150 207980 63350
rect 204150 63020 204350 63090
rect 204650 63020 204850 63090
rect 205150 63020 205350 63090
rect 205650 63020 205850 63090
rect 206150 63020 206350 63090
rect 206650 63020 206850 63090
rect 207150 63020 207350 63090
rect 207650 63020 207850 63090
rect 204150 62910 204350 62980
rect 204650 62910 204850 62980
rect 205150 62910 205350 62980
rect 205650 62910 205850 62980
rect 206150 62910 206350 62980
rect 206650 62910 206850 62980
rect 207150 62910 207350 62980
rect 207650 62910 207850 62980
rect 204020 62650 204090 62850
rect 204410 62650 204480 62850
rect 204520 62650 204590 62850
rect 204910 62650 204980 62850
rect 205020 62650 205090 62850
rect 205410 62650 205480 62850
rect 205520 62650 205590 62850
rect 205910 62650 205980 62850
rect 206020 62650 206090 62850
rect 206410 62650 206480 62850
rect 206520 62650 206590 62850
rect 206910 62650 206980 62850
rect 207020 62650 207090 62850
rect 207410 62650 207480 62850
rect 207520 62650 207590 62850
rect 207910 62650 207980 62850
rect 204150 62520 204350 62590
rect 204650 62520 204850 62590
rect 205150 62520 205350 62590
rect 205650 62520 205850 62590
rect 206150 62520 206350 62590
rect 206650 62520 206850 62590
rect 207150 62520 207350 62590
rect 207650 62520 207850 62590
rect 204150 62410 204350 62480
rect 204650 62410 204850 62480
rect 205150 62410 205350 62480
rect 205650 62410 205850 62480
rect 206150 62410 206350 62480
rect 206650 62410 206850 62480
rect 207150 62410 207350 62480
rect 207650 62410 207850 62480
rect 204020 62150 204090 62350
rect 204410 62150 204480 62350
rect 204520 62150 204590 62350
rect 204910 62150 204980 62350
rect 205020 62150 205090 62350
rect 205410 62150 205480 62350
rect 205520 62150 205590 62350
rect 205910 62150 205980 62350
rect 206020 62150 206090 62350
rect 206410 62150 206480 62350
rect 206520 62150 206590 62350
rect 206910 62150 206980 62350
rect 207020 62150 207090 62350
rect 207410 62150 207480 62350
rect 207520 62150 207590 62350
rect 207910 62150 207980 62350
rect 204150 62020 204350 62090
rect 204650 62020 204850 62090
rect 205150 62020 205350 62090
rect 205650 62020 205850 62090
rect 206150 62020 206350 62090
rect 206650 62020 206850 62090
rect 207150 62020 207350 62090
rect 207650 62020 207850 62090
rect 204150 61910 204350 61980
rect 204650 61910 204850 61980
rect 205150 61910 205350 61980
rect 205650 61910 205850 61980
rect 206150 61910 206350 61980
rect 206650 61910 206850 61980
rect 207150 61910 207350 61980
rect 207650 61910 207850 61980
rect 204020 61650 204090 61850
rect 204410 61650 204480 61850
rect 204520 61650 204590 61850
rect 204910 61650 204980 61850
rect 205020 61650 205090 61850
rect 205410 61650 205480 61850
rect 205520 61650 205590 61850
rect 205910 61650 205980 61850
rect 206020 61650 206090 61850
rect 206410 61650 206480 61850
rect 206520 61650 206590 61850
rect 206910 61650 206980 61850
rect 207020 61650 207090 61850
rect 207410 61650 207480 61850
rect 207520 61650 207590 61850
rect 207910 61650 207980 61850
rect 204150 61520 204350 61590
rect 204650 61520 204850 61590
rect 205150 61520 205350 61590
rect 205650 61520 205850 61590
rect 206150 61520 206350 61590
rect 206650 61520 206850 61590
rect 207150 61520 207350 61590
rect 207650 61520 207850 61590
rect 204150 61410 204350 61480
rect 204650 61410 204850 61480
rect 205150 61410 205350 61480
rect 205650 61410 205850 61480
rect 206150 61410 206350 61480
rect 206650 61410 206850 61480
rect 207150 61410 207350 61480
rect 207650 61410 207850 61480
rect 204020 61150 204090 61350
rect 204410 61150 204480 61350
rect 204520 61150 204590 61350
rect 204910 61150 204980 61350
rect 205020 61150 205090 61350
rect 205410 61150 205480 61350
rect 205520 61150 205590 61350
rect 205910 61150 205980 61350
rect 206020 61150 206090 61350
rect 206410 61150 206480 61350
rect 206520 61150 206590 61350
rect 206910 61150 206980 61350
rect 207020 61150 207090 61350
rect 207410 61150 207480 61350
rect 207520 61150 207590 61350
rect 207910 61150 207980 61350
rect 204150 61020 204350 61090
rect 204650 61020 204850 61090
rect 205150 61020 205350 61090
rect 205650 61020 205850 61090
rect 206150 61020 206350 61090
rect 206650 61020 206850 61090
rect 207150 61020 207350 61090
rect 207650 61020 207850 61090
rect 204150 60910 204350 60980
rect 204650 60910 204850 60980
rect 205150 60910 205350 60980
rect 205650 60910 205850 60980
rect 206150 60910 206350 60980
rect 206650 60910 206850 60980
rect 207150 60910 207350 60980
rect 207650 60910 207850 60980
rect 204020 60650 204090 60850
rect 204410 60650 204480 60850
rect 204520 60650 204590 60850
rect 204910 60650 204980 60850
rect 205020 60650 205090 60850
rect 205410 60650 205480 60850
rect 205520 60650 205590 60850
rect 205910 60650 205980 60850
rect 206020 60650 206090 60850
rect 206410 60650 206480 60850
rect 206520 60650 206590 60850
rect 206910 60650 206980 60850
rect 207020 60650 207090 60850
rect 207410 60650 207480 60850
rect 207520 60650 207590 60850
rect 207910 60650 207980 60850
rect 204150 60520 204350 60590
rect 204650 60520 204850 60590
rect 205150 60520 205350 60590
rect 205650 60520 205850 60590
rect 206150 60520 206350 60590
rect 206650 60520 206850 60590
rect 207150 60520 207350 60590
rect 207650 60520 207850 60590
rect 204150 60410 204350 60480
rect 204650 60410 204850 60480
rect 205150 60410 205350 60480
rect 205650 60410 205850 60480
rect 206150 60410 206350 60480
rect 206650 60410 206850 60480
rect 207150 60410 207350 60480
rect 207650 60410 207850 60480
rect 204020 60150 204090 60350
rect 204410 60150 204480 60350
rect 204520 60150 204590 60350
rect 204910 60150 204980 60350
rect 205020 60150 205090 60350
rect 205410 60150 205480 60350
rect 205520 60150 205590 60350
rect 205910 60150 205980 60350
rect 206020 60150 206090 60350
rect 206410 60150 206480 60350
rect 206520 60150 206590 60350
rect 206910 60150 206980 60350
rect 207020 60150 207090 60350
rect 207410 60150 207480 60350
rect 207520 60150 207590 60350
rect 207910 60150 207980 60350
rect 204150 60020 204350 60090
rect 204650 60020 204850 60090
rect 205150 60020 205350 60090
rect 205650 60020 205850 60090
rect 206150 60020 206350 60090
rect 206650 60020 206850 60090
rect 207150 60020 207350 60090
rect 207650 60020 207850 60090
rect 204150 59910 204350 59980
rect 204650 59910 204850 59980
rect 205150 59910 205350 59980
rect 205650 59910 205850 59980
rect 206150 59910 206350 59980
rect 206650 59910 206850 59980
rect 207150 59910 207350 59980
rect 207650 59910 207850 59980
rect 204020 59650 204090 59850
rect 204410 59650 204480 59850
rect 204520 59650 204590 59850
rect 204910 59650 204980 59850
rect 205020 59650 205090 59850
rect 205410 59650 205480 59850
rect 205520 59650 205590 59850
rect 205910 59650 205980 59850
rect 206020 59650 206090 59850
rect 206410 59650 206480 59850
rect 206520 59650 206590 59850
rect 206910 59650 206980 59850
rect 207020 59650 207090 59850
rect 207410 59650 207480 59850
rect 207520 59650 207590 59850
rect 207910 59650 207980 59850
rect 204150 59520 204350 59590
rect 204650 59520 204850 59590
rect 205150 59520 205350 59590
rect 205650 59520 205850 59590
rect 206150 59520 206350 59590
rect 206650 59520 206850 59590
rect 207150 59520 207350 59590
rect 207650 59520 207850 59590
rect 204150 59410 204350 59480
rect 204650 59410 204850 59480
rect 205150 59410 205350 59480
rect 205650 59410 205850 59480
rect 206150 59410 206350 59480
rect 206650 59410 206850 59480
rect 207150 59410 207350 59480
rect 207650 59410 207850 59480
rect 204020 59150 204090 59350
rect 204410 59150 204480 59350
rect 204520 59150 204590 59350
rect 204910 59150 204980 59350
rect 205020 59150 205090 59350
rect 205410 59150 205480 59350
rect 205520 59150 205590 59350
rect 205910 59150 205980 59350
rect 206020 59150 206090 59350
rect 206410 59150 206480 59350
rect 206520 59150 206590 59350
rect 206910 59150 206980 59350
rect 207020 59150 207090 59350
rect 207410 59150 207480 59350
rect 207520 59150 207590 59350
rect 207910 59150 207980 59350
rect 204150 59020 204350 59090
rect 204650 59020 204850 59090
rect 205150 59020 205350 59090
rect 205650 59020 205850 59090
rect 206150 59020 206350 59090
rect 206650 59020 206850 59090
rect 207150 59020 207350 59090
rect 207650 59020 207850 59090
rect 204150 58910 204350 58980
rect 204650 58910 204850 58980
rect 205150 58910 205350 58980
rect 205650 58910 205850 58980
rect 206150 58910 206350 58980
rect 206650 58910 206850 58980
rect 207150 58910 207350 58980
rect 207650 58910 207850 58980
rect 204020 58650 204090 58850
rect 204410 58650 204480 58850
rect 204520 58650 204590 58850
rect 204910 58650 204980 58850
rect 205020 58650 205090 58850
rect 205410 58650 205480 58850
rect 205520 58650 205590 58850
rect 205910 58650 205980 58850
rect 206020 58650 206090 58850
rect 206410 58650 206480 58850
rect 206520 58650 206590 58850
rect 206910 58650 206980 58850
rect 207020 58650 207090 58850
rect 207410 58650 207480 58850
rect 207520 58650 207590 58850
rect 207910 58650 207980 58850
rect 204150 58520 204350 58590
rect 204650 58520 204850 58590
rect 205150 58520 205350 58590
rect 205650 58520 205850 58590
rect 206150 58520 206350 58590
rect 206650 58520 206850 58590
rect 207150 58520 207350 58590
rect 207650 58520 207850 58590
rect 204150 58410 204350 58480
rect 204650 58410 204850 58480
rect 205150 58410 205350 58480
rect 205650 58410 205850 58480
rect 206150 58410 206350 58480
rect 206650 58410 206850 58480
rect 207150 58410 207350 58480
rect 207650 58410 207850 58480
rect 204020 58150 204090 58350
rect 204410 58150 204480 58350
rect 204520 58150 204590 58350
rect 204910 58150 204980 58350
rect 205020 58150 205090 58350
rect 205410 58150 205480 58350
rect 205520 58150 205590 58350
rect 205910 58150 205980 58350
rect 206020 58150 206090 58350
rect 206410 58150 206480 58350
rect 206520 58150 206590 58350
rect 206910 58150 206980 58350
rect 207020 58150 207090 58350
rect 207410 58150 207480 58350
rect 207520 58150 207590 58350
rect 207910 58150 207980 58350
rect 204150 58020 204350 58090
rect 204650 58020 204850 58090
rect 205150 58020 205350 58090
rect 205650 58020 205850 58090
rect 206150 58020 206350 58090
rect 206650 58020 206850 58090
rect 207150 58020 207350 58090
rect 207650 58020 207850 58090
rect 204150 57910 204350 57980
rect 204650 57910 204850 57980
rect 205150 57910 205350 57980
rect 205650 57910 205850 57980
rect 206150 57910 206350 57980
rect 206650 57910 206850 57980
rect 207150 57910 207350 57980
rect 207650 57910 207850 57980
rect 204020 57650 204090 57850
rect 204410 57650 204480 57850
rect 204520 57650 204590 57850
rect 204910 57650 204980 57850
rect 205020 57650 205090 57850
rect 205410 57650 205480 57850
rect 205520 57650 205590 57850
rect 205910 57650 205980 57850
rect 206020 57650 206090 57850
rect 206410 57650 206480 57850
rect 206520 57650 206590 57850
rect 206910 57650 206980 57850
rect 207020 57650 207090 57850
rect 207410 57650 207480 57850
rect 207520 57650 207590 57850
rect 207910 57650 207980 57850
rect 204150 57520 204350 57590
rect 204650 57520 204850 57590
rect 205150 57520 205350 57590
rect 205650 57520 205850 57590
rect 206150 57520 206350 57590
rect 206650 57520 206850 57590
rect 207150 57520 207350 57590
rect 207650 57520 207850 57590
rect 204150 57410 204350 57480
rect 204650 57410 204850 57480
rect 205150 57410 205350 57480
rect 205650 57410 205850 57480
rect 206150 57410 206350 57480
rect 206650 57410 206850 57480
rect 207150 57410 207350 57480
rect 207650 57410 207850 57480
rect 204020 57150 204090 57350
rect 204410 57150 204480 57350
rect 204520 57150 204590 57350
rect 204910 57150 204980 57350
rect 205020 57150 205090 57350
rect 205410 57150 205480 57350
rect 205520 57150 205590 57350
rect 205910 57150 205980 57350
rect 206020 57150 206090 57350
rect 206410 57150 206480 57350
rect 206520 57150 206590 57350
rect 206910 57150 206980 57350
rect 207020 57150 207090 57350
rect 207410 57150 207480 57350
rect 207520 57150 207590 57350
rect 207910 57150 207980 57350
rect 204150 57020 204350 57090
rect 204650 57020 204850 57090
rect 205150 57020 205350 57090
rect 205650 57020 205850 57090
rect 206150 57020 206350 57090
rect 206650 57020 206850 57090
rect 207150 57020 207350 57090
rect 207650 57020 207850 57090
rect 204150 56910 204350 56980
rect 204650 56910 204850 56980
rect 205150 56910 205350 56980
rect 205650 56910 205850 56980
rect 206150 56910 206350 56980
rect 206650 56910 206850 56980
rect 207150 56910 207350 56980
rect 207650 56910 207850 56980
rect 204020 56650 204090 56850
rect 204410 56650 204480 56850
rect 204520 56650 204590 56850
rect 204910 56650 204980 56850
rect 205020 56650 205090 56850
rect 205410 56650 205480 56850
rect 205520 56650 205590 56850
rect 205910 56650 205980 56850
rect 206020 56650 206090 56850
rect 206410 56650 206480 56850
rect 206520 56650 206590 56850
rect 206910 56650 206980 56850
rect 207020 56650 207090 56850
rect 207410 56650 207480 56850
rect 207520 56650 207590 56850
rect 207910 56650 207980 56850
rect 204150 56520 204350 56590
rect 204650 56520 204850 56590
rect 205150 56520 205350 56590
rect 205650 56520 205850 56590
rect 206150 56520 206350 56590
rect 206650 56520 206850 56590
rect 207150 56520 207350 56590
rect 207650 56520 207850 56590
rect 204150 56410 204350 56480
rect 204650 56410 204850 56480
rect 205150 56410 205350 56480
rect 205650 56410 205850 56480
rect 206150 56410 206350 56480
rect 206650 56410 206850 56480
rect 207150 56410 207350 56480
rect 207650 56410 207850 56480
rect 204020 56150 204090 56350
rect 204410 56150 204480 56350
rect 204520 56150 204590 56350
rect 204910 56150 204980 56350
rect 205020 56150 205090 56350
rect 205410 56150 205480 56350
rect 205520 56150 205590 56350
rect 205910 56150 205980 56350
rect 206020 56150 206090 56350
rect 206410 56150 206480 56350
rect 206520 56150 206590 56350
rect 206910 56150 206980 56350
rect 207020 56150 207090 56350
rect 207410 56150 207480 56350
rect 207520 56150 207590 56350
rect 207910 56150 207980 56350
rect 204150 56020 204350 56090
rect 204650 56020 204850 56090
rect 205150 56020 205350 56090
rect 205650 56020 205850 56090
rect 206150 56020 206350 56090
rect 206650 56020 206850 56090
rect 207150 56020 207350 56090
rect 207650 56020 207850 56090
rect 204150 55910 204350 55980
rect 204650 55910 204850 55980
rect 205150 55910 205350 55980
rect 205650 55910 205850 55980
rect 206150 55910 206350 55980
rect 206650 55910 206850 55980
rect 207150 55910 207350 55980
rect 207650 55910 207850 55980
rect 204020 55650 204090 55850
rect 204410 55650 204480 55850
rect 204520 55650 204590 55850
rect 204910 55650 204980 55850
rect 205020 55650 205090 55850
rect 205410 55650 205480 55850
rect 205520 55650 205590 55850
rect 205910 55650 205980 55850
rect 206020 55650 206090 55850
rect 206410 55650 206480 55850
rect 206520 55650 206590 55850
rect 206910 55650 206980 55850
rect 207020 55650 207090 55850
rect 207410 55650 207480 55850
rect 207520 55650 207590 55850
rect 207910 55650 207980 55850
rect 204150 55520 204350 55590
rect 204650 55520 204850 55590
rect 205150 55520 205350 55590
rect 205650 55520 205850 55590
rect 206150 55520 206350 55590
rect 206650 55520 206850 55590
rect 207150 55520 207350 55590
rect 207650 55520 207850 55590
rect 204150 55410 204350 55480
rect 204650 55410 204850 55480
rect 205150 55410 205350 55480
rect 205650 55410 205850 55480
rect 206150 55410 206350 55480
rect 206650 55410 206850 55480
rect 207150 55410 207350 55480
rect 207650 55410 207850 55480
rect 204020 55150 204090 55350
rect 204410 55150 204480 55350
rect 204520 55150 204590 55350
rect 204910 55150 204980 55350
rect 205020 55150 205090 55350
rect 205410 55150 205480 55350
rect 205520 55150 205590 55350
rect 205910 55150 205980 55350
rect 206020 55150 206090 55350
rect 206410 55150 206480 55350
rect 206520 55150 206590 55350
rect 206910 55150 206980 55350
rect 207020 55150 207090 55350
rect 207410 55150 207480 55350
rect 207520 55150 207590 55350
rect 207910 55150 207980 55350
rect 204150 55020 204350 55090
rect 204650 55020 204850 55090
rect 205150 55020 205350 55090
rect 205650 55020 205850 55090
rect 206150 55020 206350 55090
rect 206650 55020 206850 55090
rect 207150 55020 207350 55090
rect 207650 55020 207850 55090
rect 204150 54910 204350 54980
rect 204650 54910 204850 54980
rect 205150 54910 205350 54980
rect 205650 54910 205850 54980
rect 206150 54910 206350 54980
rect 206650 54910 206850 54980
rect 207150 54910 207350 54980
rect 207650 54910 207850 54980
rect 204020 54650 204090 54850
rect 204410 54650 204480 54850
rect 204520 54650 204590 54850
rect 204910 54650 204980 54850
rect 205020 54650 205090 54850
rect 205410 54650 205480 54850
rect 205520 54650 205590 54850
rect 205910 54650 205980 54850
rect 206020 54650 206090 54850
rect 206410 54650 206480 54850
rect 206520 54650 206590 54850
rect 206910 54650 206980 54850
rect 207020 54650 207090 54850
rect 207410 54650 207480 54850
rect 207520 54650 207590 54850
rect 207910 54650 207980 54850
rect 204150 54520 204350 54590
rect 204650 54520 204850 54590
rect 205150 54520 205350 54590
rect 205650 54520 205850 54590
rect 206150 54520 206350 54590
rect 206650 54520 206850 54590
rect 207150 54520 207350 54590
rect 207650 54520 207850 54590
rect 204150 54410 204350 54480
rect 204650 54410 204850 54480
rect 205150 54410 205350 54480
rect 205650 54410 205850 54480
rect 206150 54410 206350 54480
rect 206650 54410 206850 54480
rect 207150 54410 207350 54480
rect 207650 54410 207850 54480
rect 204020 54150 204090 54350
rect 204410 54150 204480 54350
rect 204520 54150 204590 54350
rect 204910 54150 204980 54350
rect 205020 54150 205090 54350
rect 205410 54150 205480 54350
rect 205520 54150 205590 54350
rect 205910 54150 205980 54350
rect 206020 54150 206090 54350
rect 206410 54150 206480 54350
rect 206520 54150 206590 54350
rect 206910 54150 206980 54350
rect 207020 54150 207090 54350
rect 207410 54150 207480 54350
rect 207520 54150 207590 54350
rect 207910 54150 207980 54350
rect 204150 54020 204350 54090
rect 204650 54020 204850 54090
rect 205150 54020 205350 54090
rect 205650 54020 205850 54090
rect 206150 54020 206350 54090
rect 206650 54020 206850 54090
rect 207150 54020 207350 54090
rect 207650 54020 207850 54090
rect 204150 53910 204350 53980
rect 204650 53910 204850 53980
rect 205150 53910 205350 53980
rect 205650 53910 205850 53980
rect 206150 53910 206350 53980
rect 206650 53910 206850 53980
rect 207150 53910 207350 53980
rect 207650 53910 207850 53980
rect 204020 53650 204090 53850
rect 204410 53650 204480 53850
rect 204520 53650 204590 53850
rect 204910 53650 204980 53850
rect 205020 53650 205090 53850
rect 205410 53650 205480 53850
rect 205520 53650 205590 53850
rect 205910 53650 205980 53850
rect 206020 53650 206090 53850
rect 206410 53650 206480 53850
rect 206520 53650 206590 53850
rect 206910 53650 206980 53850
rect 207020 53650 207090 53850
rect 207410 53650 207480 53850
rect 207520 53650 207590 53850
rect 207910 53650 207980 53850
rect 204150 53520 204350 53590
rect 204650 53520 204850 53590
rect 205150 53520 205350 53590
rect 205650 53520 205850 53590
rect 206150 53520 206350 53590
rect 206650 53520 206850 53590
rect 207150 53520 207350 53590
rect 207650 53520 207850 53590
rect 204150 53410 204350 53480
rect 204650 53410 204850 53480
rect 205150 53410 205350 53480
rect 205650 53410 205850 53480
rect 206150 53410 206350 53480
rect 206650 53410 206850 53480
rect 207150 53410 207350 53480
rect 207650 53410 207850 53480
rect 204020 53150 204090 53350
rect 204410 53150 204480 53350
rect 204520 53150 204590 53350
rect 204910 53150 204980 53350
rect 205020 53150 205090 53350
rect 205410 53150 205480 53350
rect 205520 53150 205590 53350
rect 205910 53150 205980 53350
rect 206020 53150 206090 53350
rect 206410 53150 206480 53350
rect 206520 53150 206590 53350
rect 206910 53150 206980 53350
rect 207020 53150 207090 53350
rect 207410 53150 207480 53350
rect 207520 53150 207590 53350
rect 207910 53150 207980 53350
rect 204150 53020 204350 53090
rect 204650 53020 204850 53090
rect 205150 53020 205350 53090
rect 205650 53020 205850 53090
rect 206150 53020 206350 53090
rect 206650 53020 206850 53090
rect 207150 53020 207350 53090
rect 207650 53020 207850 53090
rect 204150 52910 204350 52980
rect 204650 52910 204850 52980
rect 205150 52910 205350 52980
rect 205650 52910 205850 52980
rect 206150 52910 206350 52980
rect 206650 52910 206850 52980
rect 207150 52910 207350 52980
rect 207650 52910 207850 52980
rect 204020 52650 204090 52850
rect 204410 52650 204480 52850
rect 204520 52650 204590 52850
rect 204910 52650 204980 52850
rect 205020 52650 205090 52850
rect 205410 52650 205480 52850
rect 205520 52650 205590 52850
rect 205910 52650 205980 52850
rect 206020 52650 206090 52850
rect 206410 52650 206480 52850
rect 206520 52650 206590 52850
rect 206910 52650 206980 52850
rect 207020 52650 207090 52850
rect 207410 52650 207480 52850
rect 207520 52650 207590 52850
rect 207910 52650 207980 52850
rect 204150 52520 204350 52590
rect 204650 52520 204850 52590
rect 205150 52520 205350 52590
rect 205650 52520 205850 52590
rect 206150 52520 206350 52590
rect 206650 52520 206850 52590
rect 207150 52520 207350 52590
rect 207650 52520 207850 52590
rect 204150 52410 204350 52480
rect 204650 52410 204850 52480
rect 205150 52410 205350 52480
rect 205650 52410 205850 52480
rect 206150 52410 206350 52480
rect 206650 52410 206850 52480
rect 207150 52410 207350 52480
rect 207650 52410 207850 52480
rect 204020 52150 204090 52350
rect 204410 52150 204480 52350
rect 204520 52150 204590 52350
rect 204910 52150 204980 52350
rect 205020 52150 205090 52350
rect 205410 52150 205480 52350
rect 205520 52150 205590 52350
rect 205910 52150 205980 52350
rect 206020 52150 206090 52350
rect 206410 52150 206480 52350
rect 206520 52150 206590 52350
rect 206910 52150 206980 52350
rect 207020 52150 207090 52350
rect 207410 52150 207480 52350
rect 207520 52150 207590 52350
rect 207910 52150 207980 52350
rect 204150 52020 204350 52090
rect 204650 52020 204850 52090
rect 205150 52020 205350 52090
rect 205650 52020 205850 52090
rect 206150 52020 206350 52090
rect 206650 52020 206850 52090
rect 207150 52020 207350 52090
rect 207650 52020 207850 52090
rect 204150 51910 204350 51980
rect 204650 51910 204850 51980
rect 205150 51910 205350 51980
rect 205650 51910 205850 51980
rect 206150 51910 206350 51980
rect 206650 51910 206850 51980
rect 207150 51910 207350 51980
rect 207650 51910 207850 51980
rect 204020 51650 204090 51850
rect 204410 51650 204480 51850
rect 204520 51650 204590 51850
rect 204910 51650 204980 51850
rect 205020 51650 205090 51850
rect 205410 51650 205480 51850
rect 205520 51650 205590 51850
rect 205910 51650 205980 51850
rect 206020 51650 206090 51850
rect 206410 51650 206480 51850
rect 206520 51650 206590 51850
rect 206910 51650 206980 51850
rect 207020 51650 207090 51850
rect 207410 51650 207480 51850
rect 207520 51650 207590 51850
rect 207910 51650 207980 51850
rect 204150 51520 204350 51590
rect 204650 51520 204850 51590
rect 205150 51520 205350 51590
rect 205650 51520 205850 51590
rect 206150 51520 206350 51590
rect 206650 51520 206850 51590
rect 207150 51520 207350 51590
rect 207650 51520 207850 51590
rect 204150 51410 204350 51480
rect 204650 51410 204850 51480
rect 205150 51410 205350 51480
rect 205650 51410 205850 51480
rect 206150 51410 206350 51480
rect 206650 51410 206850 51480
rect 207150 51410 207350 51480
rect 207650 51410 207850 51480
rect 204020 51150 204090 51350
rect 204410 51150 204480 51350
rect 204520 51150 204590 51350
rect 204910 51150 204980 51350
rect 205020 51150 205090 51350
rect 205410 51150 205480 51350
rect 205520 51150 205590 51350
rect 205910 51150 205980 51350
rect 206020 51150 206090 51350
rect 206410 51150 206480 51350
rect 206520 51150 206590 51350
rect 206910 51150 206980 51350
rect 207020 51150 207090 51350
rect 207410 51150 207480 51350
rect 207520 51150 207590 51350
rect 207910 51150 207980 51350
rect 204150 51020 204350 51090
rect 204650 51020 204850 51090
rect 205150 51020 205350 51090
rect 205650 51020 205850 51090
rect 206150 51020 206350 51090
rect 206650 51020 206850 51090
rect 207150 51020 207350 51090
rect 207650 51020 207850 51090
rect 204150 50910 204350 50980
rect 204650 50910 204850 50980
rect 205150 50910 205350 50980
rect 205650 50910 205850 50980
rect 206150 50910 206350 50980
rect 206650 50910 206850 50980
rect 207150 50910 207350 50980
rect 207650 50910 207850 50980
rect 204020 50650 204090 50850
rect 204410 50650 204480 50850
rect 204520 50650 204590 50850
rect 204910 50650 204980 50850
rect 205020 50650 205090 50850
rect 205410 50650 205480 50850
rect 205520 50650 205590 50850
rect 205910 50650 205980 50850
rect 206020 50650 206090 50850
rect 206410 50650 206480 50850
rect 206520 50650 206590 50850
rect 206910 50650 206980 50850
rect 207020 50650 207090 50850
rect 207410 50650 207480 50850
rect 207520 50650 207590 50850
rect 207910 50650 207980 50850
rect 204150 50520 204350 50590
rect 204650 50520 204850 50590
rect 205150 50520 205350 50590
rect 205650 50520 205850 50590
rect 206150 50520 206350 50590
rect 206650 50520 206850 50590
rect 207150 50520 207350 50590
rect 207650 50520 207850 50590
rect 204150 50410 204350 50480
rect 204650 50410 204850 50480
rect 205150 50410 205350 50480
rect 205650 50410 205850 50480
rect 206150 50410 206350 50480
rect 206650 50410 206850 50480
rect 207150 50410 207350 50480
rect 207650 50410 207850 50480
rect 204020 50150 204090 50350
rect 204410 50150 204480 50350
rect 204520 50150 204590 50350
rect 204910 50150 204980 50350
rect 205020 50150 205090 50350
rect 205410 50150 205480 50350
rect 205520 50150 205590 50350
rect 205910 50150 205980 50350
rect 206020 50150 206090 50350
rect 206410 50150 206480 50350
rect 206520 50150 206590 50350
rect 206910 50150 206980 50350
rect 207020 50150 207090 50350
rect 207410 50150 207480 50350
rect 207520 50150 207590 50350
rect 207910 50150 207980 50350
rect 204150 50020 204350 50090
rect 204650 50020 204850 50090
rect 205150 50020 205350 50090
rect 205650 50020 205850 50090
rect 206150 50020 206350 50090
rect 206650 50020 206850 50090
rect 207150 50020 207350 50090
rect 207650 50020 207850 50090
rect 204150 49910 204350 49980
rect 204650 49910 204850 49980
rect 205150 49910 205350 49980
rect 205650 49910 205850 49980
rect 206150 49910 206350 49980
rect 206650 49910 206850 49980
rect 207150 49910 207350 49980
rect 207650 49910 207850 49980
rect 204020 49650 204090 49850
rect 204410 49650 204480 49850
rect 204520 49650 204590 49850
rect 204910 49650 204980 49850
rect 205020 49650 205090 49850
rect 205410 49650 205480 49850
rect 205520 49650 205590 49850
rect 205910 49650 205980 49850
rect 206020 49650 206090 49850
rect 206410 49650 206480 49850
rect 206520 49650 206590 49850
rect 206910 49650 206980 49850
rect 207020 49650 207090 49850
rect 207410 49650 207480 49850
rect 207520 49650 207590 49850
rect 207910 49650 207980 49850
rect 204150 49520 204350 49590
rect 204650 49520 204850 49590
rect 205150 49520 205350 49590
rect 205650 49520 205850 49590
rect 206150 49520 206350 49590
rect 206650 49520 206850 49590
rect 207150 49520 207350 49590
rect 207650 49520 207850 49590
rect 204150 49410 204350 49480
rect 204650 49410 204850 49480
rect 205150 49410 205350 49480
rect 205650 49410 205850 49480
rect 206150 49410 206350 49480
rect 206650 49410 206850 49480
rect 207150 49410 207350 49480
rect 207650 49410 207850 49480
rect 204020 49150 204090 49350
rect 204410 49150 204480 49350
rect 204520 49150 204590 49350
rect 204910 49150 204980 49350
rect 205020 49150 205090 49350
rect 205410 49150 205480 49350
rect 205520 49150 205590 49350
rect 205910 49150 205980 49350
rect 206020 49150 206090 49350
rect 206410 49150 206480 49350
rect 206520 49150 206590 49350
rect 206910 49150 206980 49350
rect 207020 49150 207090 49350
rect 207410 49150 207480 49350
rect 207520 49150 207590 49350
rect 207910 49150 207980 49350
rect 204150 49020 204350 49090
rect 204650 49020 204850 49090
rect 205150 49020 205350 49090
rect 205650 49020 205850 49090
rect 206150 49020 206350 49090
rect 206650 49020 206850 49090
rect 207150 49020 207350 49090
rect 207650 49020 207850 49090
rect 204150 48910 204350 48980
rect 204650 48910 204850 48980
rect 205150 48910 205350 48980
rect 205650 48910 205850 48980
rect 206150 48910 206350 48980
rect 206650 48910 206850 48980
rect 207150 48910 207350 48980
rect 207650 48910 207850 48980
rect 204020 48650 204090 48850
rect 204410 48650 204480 48850
rect 204520 48650 204590 48850
rect 204910 48650 204980 48850
rect 205020 48650 205090 48850
rect 205410 48650 205480 48850
rect 205520 48650 205590 48850
rect 205910 48650 205980 48850
rect 206020 48650 206090 48850
rect 206410 48650 206480 48850
rect 206520 48650 206590 48850
rect 206910 48650 206980 48850
rect 207020 48650 207090 48850
rect 207410 48650 207480 48850
rect 207520 48650 207590 48850
rect 207910 48650 207980 48850
rect 204150 48520 204350 48590
rect 204650 48520 204850 48590
rect 205150 48520 205350 48590
rect 205650 48520 205850 48590
rect 206150 48520 206350 48590
rect 206650 48520 206850 48590
rect 207150 48520 207350 48590
rect 207650 48520 207850 48590
rect 204150 48410 204350 48480
rect 204650 48410 204850 48480
rect 205150 48410 205350 48480
rect 205650 48410 205850 48480
rect 206150 48410 206350 48480
rect 206650 48410 206850 48480
rect 207150 48410 207350 48480
rect 207650 48410 207850 48480
rect 204020 48150 204090 48350
rect 204410 48150 204480 48350
rect 204520 48150 204590 48350
rect 204910 48150 204980 48350
rect 205020 48150 205090 48350
rect 205410 48150 205480 48350
rect 205520 48150 205590 48350
rect 205910 48150 205980 48350
rect 206020 48150 206090 48350
rect 206410 48150 206480 48350
rect 206520 48150 206590 48350
rect 206910 48150 206980 48350
rect 207020 48150 207090 48350
rect 207410 48150 207480 48350
rect 207520 48150 207590 48350
rect 207910 48150 207980 48350
rect 204150 48020 204350 48090
rect 204650 48020 204850 48090
rect 205150 48020 205350 48090
rect 205650 48020 205850 48090
rect 206150 48020 206350 48090
rect 206650 48020 206850 48090
rect 207150 48020 207350 48090
rect 207650 48020 207850 48090
rect 204150 47910 204350 47980
rect 204650 47910 204850 47980
rect 205150 47910 205350 47980
rect 205650 47910 205850 47980
rect 206150 47910 206350 47980
rect 206650 47910 206850 47980
rect 207150 47910 207350 47980
rect 207650 47910 207850 47980
rect 204020 47650 204090 47850
rect 204410 47650 204480 47850
rect 204520 47650 204590 47850
rect 204910 47650 204980 47850
rect 205020 47650 205090 47850
rect 205410 47650 205480 47850
rect 205520 47650 205590 47850
rect 205910 47650 205980 47850
rect 206020 47650 206090 47850
rect 206410 47650 206480 47850
rect 206520 47650 206590 47850
rect 206910 47650 206980 47850
rect 207020 47650 207090 47850
rect 207410 47650 207480 47850
rect 207520 47650 207590 47850
rect 207910 47650 207980 47850
rect 204150 47520 204350 47590
rect 204650 47520 204850 47590
rect 205150 47520 205350 47590
rect 205650 47520 205850 47590
rect 206150 47520 206350 47590
rect 206650 47520 206850 47590
rect 207150 47520 207350 47590
rect 207650 47520 207850 47590
rect 204150 47410 204350 47480
rect 204650 47410 204850 47480
rect 205150 47410 205350 47480
rect 205650 47410 205850 47480
rect 206150 47410 206350 47480
rect 206650 47410 206850 47480
rect 207150 47410 207350 47480
rect 207650 47410 207850 47480
rect 204020 47150 204090 47350
rect 204410 47150 204480 47350
rect 204520 47150 204590 47350
rect 204910 47150 204980 47350
rect 205020 47150 205090 47350
rect 205410 47150 205480 47350
rect 205520 47150 205590 47350
rect 205910 47150 205980 47350
rect 206020 47150 206090 47350
rect 206410 47150 206480 47350
rect 206520 47150 206590 47350
rect 206910 47150 206980 47350
rect 207020 47150 207090 47350
rect 207410 47150 207480 47350
rect 207520 47150 207590 47350
rect 207910 47150 207980 47350
rect 204150 47020 204350 47090
rect 204650 47020 204850 47090
rect 205150 47020 205350 47090
rect 205650 47020 205850 47090
rect 206150 47020 206350 47090
rect 206650 47020 206850 47090
rect 207150 47020 207350 47090
rect 207650 47020 207850 47090
rect 204150 46910 204350 46980
rect 204650 46910 204850 46980
rect 205150 46910 205350 46980
rect 205650 46910 205850 46980
rect 206150 46910 206350 46980
rect 206650 46910 206850 46980
rect 207150 46910 207350 46980
rect 207650 46910 207850 46980
rect 204020 46650 204090 46850
rect 204410 46650 204480 46850
rect 204520 46650 204590 46850
rect 204910 46650 204980 46850
rect 205020 46650 205090 46850
rect 205410 46650 205480 46850
rect 205520 46650 205590 46850
rect 205910 46650 205980 46850
rect 206020 46650 206090 46850
rect 206410 46650 206480 46850
rect 206520 46650 206590 46850
rect 206910 46650 206980 46850
rect 207020 46650 207090 46850
rect 207410 46650 207480 46850
rect 207520 46650 207590 46850
rect 207910 46650 207980 46850
rect 204150 46520 204350 46590
rect 204650 46520 204850 46590
rect 205150 46520 205350 46590
rect 205650 46520 205850 46590
rect 206150 46520 206350 46590
rect 206650 46520 206850 46590
rect 207150 46520 207350 46590
rect 207650 46520 207850 46590
rect 204150 46410 204350 46480
rect 204650 46410 204850 46480
rect 205150 46410 205350 46480
rect 205650 46410 205850 46480
rect 206150 46410 206350 46480
rect 206650 46410 206850 46480
rect 207150 46410 207350 46480
rect 207650 46410 207850 46480
rect 204020 46150 204090 46350
rect 204410 46150 204480 46350
rect 204520 46150 204590 46350
rect 204910 46150 204980 46350
rect 205020 46150 205090 46350
rect 205410 46150 205480 46350
rect 205520 46150 205590 46350
rect 205910 46150 205980 46350
rect 206020 46150 206090 46350
rect 206410 46150 206480 46350
rect 206520 46150 206590 46350
rect 206910 46150 206980 46350
rect 207020 46150 207090 46350
rect 207410 46150 207480 46350
rect 207520 46150 207590 46350
rect 207910 46150 207980 46350
rect 204150 46020 204350 46090
rect 204650 46020 204850 46090
rect 205150 46020 205350 46090
rect 205650 46020 205850 46090
rect 206150 46020 206350 46090
rect 206650 46020 206850 46090
rect 207150 46020 207350 46090
rect 207650 46020 207850 46090
rect 204150 45910 204350 45980
rect 204650 45910 204850 45980
rect 205150 45910 205350 45980
rect 205650 45910 205850 45980
rect 206150 45910 206350 45980
rect 206650 45910 206850 45980
rect 207150 45910 207350 45980
rect 207650 45910 207850 45980
rect 204020 45650 204090 45850
rect 204410 45650 204480 45850
rect 204520 45650 204590 45850
rect 204910 45650 204980 45850
rect 205020 45650 205090 45850
rect 205410 45650 205480 45850
rect 205520 45650 205590 45850
rect 205910 45650 205980 45850
rect 206020 45650 206090 45850
rect 206410 45650 206480 45850
rect 206520 45650 206590 45850
rect 206910 45650 206980 45850
rect 207020 45650 207090 45850
rect 207410 45650 207480 45850
rect 207520 45650 207590 45850
rect 207910 45650 207980 45850
rect 204150 45520 204350 45590
rect 204650 45520 204850 45590
rect 205150 45520 205350 45590
rect 205650 45520 205850 45590
rect 206150 45520 206350 45590
rect 206650 45520 206850 45590
rect 207150 45520 207350 45590
rect 207650 45520 207850 45590
rect 204150 45410 204350 45480
rect 204650 45410 204850 45480
rect 205150 45410 205350 45480
rect 205650 45410 205850 45480
rect 206150 45410 206350 45480
rect 206650 45410 206850 45480
rect 207150 45410 207350 45480
rect 207650 45410 207850 45480
rect 204020 45150 204090 45350
rect 204410 45150 204480 45350
rect 204520 45150 204590 45350
rect 204910 45150 204980 45350
rect 205020 45150 205090 45350
rect 205410 45150 205480 45350
rect 205520 45150 205590 45350
rect 205910 45150 205980 45350
rect 206020 45150 206090 45350
rect 206410 45150 206480 45350
rect 206520 45150 206590 45350
rect 206910 45150 206980 45350
rect 207020 45150 207090 45350
rect 207410 45150 207480 45350
rect 207520 45150 207590 45350
rect 207910 45150 207980 45350
rect 204150 45020 204350 45090
rect 204650 45020 204850 45090
rect 205150 45020 205350 45090
rect 205650 45020 205850 45090
rect 206150 45020 206350 45090
rect 206650 45020 206850 45090
rect 207150 45020 207350 45090
rect 207650 45020 207850 45090
rect 204150 44910 204350 44980
rect 204650 44910 204850 44980
rect 205150 44910 205350 44980
rect 205650 44910 205850 44980
rect 206150 44910 206350 44980
rect 206650 44910 206850 44980
rect 207150 44910 207350 44980
rect 207650 44910 207850 44980
rect 204020 44650 204090 44850
rect 204410 44650 204480 44850
rect 204520 44650 204590 44850
rect 204910 44650 204980 44850
rect 205020 44650 205090 44850
rect 205410 44650 205480 44850
rect 205520 44650 205590 44850
rect 205910 44650 205980 44850
rect 206020 44650 206090 44850
rect 206410 44650 206480 44850
rect 206520 44650 206590 44850
rect 206910 44650 206980 44850
rect 207020 44650 207090 44850
rect 207410 44650 207480 44850
rect 207520 44650 207590 44850
rect 207910 44650 207980 44850
rect 204150 44520 204350 44590
rect 204650 44520 204850 44590
rect 205150 44520 205350 44590
rect 205650 44520 205850 44590
rect 206150 44520 206350 44590
rect 206650 44520 206850 44590
rect 207150 44520 207350 44590
rect 207650 44520 207850 44590
rect 204150 44410 204350 44480
rect 204650 44410 204850 44480
rect 205150 44410 205350 44480
rect 205650 44410 205850 44480
rect 206150 44410 206350 44480
rect 206650 44410 206850 44480
rect 207150 44410 207350 44480
rect 207650 44410 207850 44480
rect 204020 44150 204090 44350
rect 204410 44150 204480 44350
rect 204520 44150 204590 44350
rect 204910 44150 204980 44350
rect 205020 44150 205090 44350
rect 205410 44150 205480 44350
rect 205520 44150 205590 44350
rect 205910 44150 205980 44350
rect 206020 44150 206090 44350
rect 206410 44150 206480 44350
rect 206520 44150 206590 44350
rect 206910 44150 206980 44350
rect 207020 44150 207090 44350
rect 207410 44150 207480 44350
rect 207520 44150 207590 44350
rect 207910 44150 207980 44350
rect 204150 44020 204350 44090
rect 204650 44020 204850 44090
rect 205150 44020 205350 44090
rect 205650 44020 205850 44090
rect 206150 44020 206350 44090
rect 206650 44020 206850 44090
rect 207150 44020 207350 44090
rect 207650 44020 207850 44090
rect 204150 43910 204350 43980
rect 204650 43910 204850 43980
rect 205150 43910 205350 43980
rect 205650 43910 205850 43980
rect 206150 43910 206350 43980
rect 206650 43910 206850 43980
rect 207150 43910 207350 43980
rect 207650 43910 207850 43980
rect 204020 43650 204090 43850
rect 204410 43650 204480 43850
rect 204520 43650 204590 43850
rect 204910 43650 204980 43850
rect 205020 43650 205090 43850
rect 205410 43650 205480 43850
rect 205520 43650 205590 43850
rect 205910 43650 205980 43850
rect 206020 43650 206090 43850
rect 206410 43650 206480 43850
rect 206520 43650 206590 43850
rect 206910 43650 206980 43850
rect 207020 43650 207090 43850
rect 207410 43650 207480 43850
rect 207520 43650 207590 43850
rect 207910 43650 207980 43850
rect 204150 43520 204350 43590
rect 204650 43520 204850 43590
rect 205150 43520 205350 43590
rect 205650 43520 205850 43590
rect 206150 43520 206350 43590
rect 206650 43520 206850 43590
rect 207150 43520 207350 43590
rect 207650 43520 207850 43590
rect 204150 43410 204350 43480
rect 204650 43410 204850 43480
rect 205150 43410 205350 43480
rect 205650 43410 205850 43480
rect 206150 43410 206350 43480
rect 206650 43410 206850 43480
rect 207150 43410 207350 43480
rect 207650 43410 207850 43480
rect 204020 43150 204090 43350
rect 204410 43150 204480 43350
rect 204520 43150 204590 43350
rect 204910 43150 204980 43350
rect 205020 43150 205090 43350
rect 205410 43150 205480 43350
rect 205520 43150 205590 43350
rect 205910 43150 205980 43350
rect 206020 43150 206090 43350
rect 206410 43150 206480 43350
rect 206520 43150 206590 43350
rect 206910 43150 206980 43350
rect 207020 43150 207090 43350
rect 207410 43150 207480 43350
rect 207520 43150 207590 43350
rect 207910 43150 207980 43350
rect 204150 43020 204350 43090
rect 204650 43020 204850 43090
rect 205150 43020 205350 43090
rect 205650 43020 205850 43090
rect 206150 43020 206350 43090
rect 206650 43020 206850 43090
rect 207150 43020 207350 43090
rect 207650 43020 207850 43090
rect 204150 42910 204350 42980
rect 204650 42910 204850 42980
rect 205150 42910 205350 42980
rect 205650 42910 205850 42980
rect 206150 42910 206350 42980
rect 206650 42910 206850 42980
rect 207150 42910 207350 42980
rect 207650 42910 207850 42980
rect 204020 42650 204090 42850
rect 204410 42650 204480 42850
rect 204520 42650 204590 42850
rect 204910 42650 204980 42850
rect 205020 42650 205090 42850
rect 205410 42650 205480 42850
rect 205520 42650 205590 42850
rect 205910 42650 205980 42850
rect 206020 42650 206090 42850
rect 206410 42650 206480 42850
rect 206520 42650 206590 42850
rect 206910 42650 206980 42850
rect 207020 42650 207090 42850
rect 207410 42650 207480 42850
rect 207520 42650 207590 42850
rect 207910 42650 207980 42850
rect 204150 42520 204350 42590
rect 204650 42520 204850 42590
rect 205150 42520 205350 42590
rect 205650 42520 205850 42590
rect 206150 42520 206350 42590
rect 206650 42520 206850 42590
rect 207150 42520 207350 42590
rect 207650 42520 207850 42590
rect 204150 42410 204350 42480
rect 204650 42410 204850 42480
rect 205150 42410 205350 42480
rect 205650 42410 205850 42480
rect 206150 42410 206350 42480
rect 206650 42410 206850 42480
rect 207150 42410 207350 42480
rect 207650 42410 207850 42480
rect 204020 42150 204090 42350
rect 204410 42150 204480 42350
rect 204520 42150 204590 42350
rect 204910 42150 204980 42350
rect 205020 42150 205090 42350
rect 205410 42150 205480 42350
rect 205520 42150 205590 42350
rect 205910 42150 205980 42350
rect 206020 42150 206090 42350
rect 206410 42150 206480 42350
rect 206520 42150 206590 42350
rect 206910 42150 206980 42350
rect 207020 42150 207090 42350
rect 207410 42150 207480 42350
rect 207520 42150 207590 42350
rect 207910 42150 207980 42350
rect 204150 42020 204350 42090
rect 204650 42020 204850 42090
rect 205150 42020 205350 42090
rect 205650 42020 205850 42090
rect 206150 42020 206350 42090
rect 206650 42020 206850 42090
rect 207150 42020 207350 42090
rect 207650 42020 207850 42090
rect 204150 41910 204350 41980
rect 204650 41910 204850 41980
rect 205150 41910 205350 41980
rect 205650 41910 205850 41980
rect 206150 41910 206350 41980
rect 206650 41910 206850 41980
rect 207150 41910 207350 41980
rect 207650 41910 207850 41980
rect 204020 41650 204090 41850
rect 204410 41650 204480 41850
rect 204520 41650 204590 41850
rect 204910 41650 204980 41850
rect 205020 41650 205090 41850
rect 205410 41650 205480 41850
rect 205520 41650 205590 41850
rect 205910 41650 205980 41850
rect 206020 41650 206090 41850
rect 206410 41650 206480 41850
rect 206520 41650 206590 41850
rect 206910 41650 206980 41850
rect 207020 41650 207090 41850
rect 207410 41650 207480 41850
rect 207520 41650 207590 41850
rect 207910 41650 207980 41850
rect 204150 41520 204350 41590
rect 204650 41520 204850 41590
rect 205150 41520 205350 41590
rect 205650 41520 205850 41590
rect 206150 41520 206350 41590
rect 206650 41520 206850 41590
rect 207150 41520 207350 41590
rect 207650 41520 207850 41590
rect 204150 41410 204350 41480
rect 204650 41410 204850 41480
rect 205150 41410 205350 41480
rect 205650 41410 205850 41480
rect 206150 41410 206350 41480
rect 206650 41410 206850 41480
rect 207150 41410 207350 41480
rect 207650 41410 207850 41480
rect 204020 41150 204090 41350
rect 204410 41150 204480 41350
rect 204520 41150 204590 41350
rect 204910 41150 204980 41350
rect 205020 41150 205090 41350
rect 205410 41150 205480 41350
rect 205520 41150 205590 41350
rect 205910 41150 205980 41350
rect 206020 41150 206090 41350
rect 206410 41150 206480 41350
rect 206520 41150 206590 41350
rect 206910 41150 206980 41350
rect 207020 41150 207090 41350
rect 207410 41150 207480 41350
rect 207520 41150 207590 41350
rect 207910 41150 207980 41350
rect 204150 41020 204350 41090
rect 204650 41020 204850 41090
rect 205150 41020 205350 41090
rect 205650 41020 205850 41090
rect 206150 41020 206350 41090
rect 206650 41020 206850 41090
rect 207150 41020 207350 41090
rect 207650 41020 207850 41090
rect 204150 40910 204350 40980
rect 204650 40910 204850 40980
rect 205150 40910 205350 40980
rect 205650 40910 205850 40980
rect 206150 40910 206350 40980
rect 206650 40910 206850 40980
rect 207150 40910 207350 40980
rect 207650 40910 207850 40980
rect 204020 40650 204090 40850
rect 204410 40650 204480 40850
rect 204520 40650 204590 40850
rect 204910 40650 204980 40850
rect 205020 40650 205090 40850
rect 205410 40650 205480 40850
rect 205520 40650 205590 40850
rect 205910 40650 205980 40850
rect 206020 40650 206090 40850
rect 206410 40650 206480 40850
rect 206520 40650 206590 40850
rect 206910 40650 206980 40850
rect 207020 40650 207090 40850
rect 207410 40650 207480 40850
rect 207520 40650 207590 40850
rect 207910 40650 207980 40850
rect 204150 40520 204350 40590
rect 204650 40520 204850 40590
rect 205150 40520 205350 40590
rect 205650 40520 205850 40590
rect 206150 40520 206350 40590
rect 206650 40520 206850 40590
rect 207150 40520 207350 40590
rect 207650 40520 207850 40590
rect 204150 40410 204350 40480
rect 204650 40410 204850 40480
rect 205150 40410 205350 40480
rect 205650 40410 205850 40480
rect 206150 40410 206350 40480
rect 206650 40410 206850 40480
rect 207150 40410 207350 40480
rect 207650 40410 207850 40480
rect 204020 40150 204090 40350
rect 204410 40150 204480 40350
rect 204520 40150 204590 40350
rect 204910 40150 204980 40350
rect 205020 40150 205090 40350
rect 205410 40150 205480 40350
rect 205520 40150 205590 40350
rect 205910 40150 205980 40350
rect 206020 40150 206090 40350
rect 206410 40150 206480 40350
rect 206520 40150 206590 40350
rect 206910 40150 206980 40350
rect 207020 40150 207090 40350
rect 207410 40150 207480 40350
rect 207520 40150 207590 40350
rect 207910 40150 207980 40350
rect 204150 40020 204350 40090
rect 204650 40020 204850 40090
rect 205150 40020 205350 40090
rect 205650 40020 205850 40090
rect 206150 40020 206350 40090
rect 206650 40020 206850 40090
rect 207150 40020 207350 40090
rect 207650 40020 207850 40090
rect 204150 39910 204350 39980
rect 204650 39910 204850 39980
rect 205150 39910 205350 39980
rect 205650 39910 205850 39980
rect 206150 39910 206350 39980
rect 206650 39910 206850 39980
rect 207150 39910 207350 39980
rect 207650 39910 207850 39980
rect 204020 39650 204090 39850
rect 204410 39650 204480 39850
rect 204520 39650 204590 39850
rect 204910 39650 204980 39850
rect 205020 39650 205090 39850
rect 205410 39650 205480 39850
rect 205520 39650 205590 39850
rect 205910 39650 205980 39850
rect 206020 39650 206090 39850
rect 206410 39650 206480 39850
rect 206520 39650 206590 39850
rect 206910 39650 206980 39850
rect 207020 39650 207090 39850
rect 207410 39650 207480 39850
rect 207520 39650 207590 39850
rect 207910 39650 207980 39850
rect 204150 39520 204350 39590
rect 204650 39520 204850 39590
rect 205150 39520 205350 39590
rect 205650 39520 205850 39590
rect 206150 39520 206350 39590
rect 206650 39520 206850 39590
rect 207150 39520 207350 39590
rect 207650 39520 207850 39590
rect 204150 39410 204350 39480
rect 204650 39410 204850 39480
rect 205150 39410 205350 39480
rect 205650 39410 205850 39480
rect 206150 39410 206350 39480
rect 206650 39410 206850 39480
rect 207150 39410 207350 39480
rect 207650 39410 207850 39480
rect 204020 39150 204090 39350
rect 204410 39150 204480 39350
rect 204520 39150 204590 39350
rect 204910 39150 204980 39350
rect 205020 39150 205090 39350
rect 205410 39150 205480 39350
rect 205520 39150 205590 39350
rect 205910 39150 205980 39350
rect 206020 39150 206090 39350
rect 206410 39150 206480 39350
rect 206520 39150 206590 39350
rect 206910 39150 206980 39350
rect 207020 39150 207090 39350
rect 207410 39150 207480 39350
rect 207520 39150 207590 39350
rect 207910 39150 207980 39350
rect 204150 39020 204350 39090
rect 204650 39020 204850 39090
rect 205150 39020 205350 39090
rect 205650 39020 205850 39090
rect 206150 39020 206350 39090
rect 206650 39020 206850 39090
rect 207150 39020 207350 39090
rect 207650 39020 207850 39090
rect 204150 38910 204350 38980
rect 204650 38910 204850 38980
rect 205150 38910 205350 38980
rect 205650 38910 205850 38980
rect 206150 38910 206350 38980
rect 206650 38910 206850 38980
rect 207150 38910 207350 38980
rect 207650 38910 207850 38980
rect 204020 38650 204090 38850
rect 204410 38650 204480 38850
rect 204520 38650 204590 38850
rect 204910 38650 204980 38850
rect 205020 38650 205090 38850
rect 205410 38650 205480 38850
rect 205520 38650 205590 38850
rect 205910 38650 205980 38850
rect 206020 38650 206090 38850
rect 206410 38650 206480 38850
rect 206520 38650 206590 38850
rect 206910 38650 206980 38850
rect 207020 38650 207090 38850
rect 207410 38650 207480 38850
rect 207520 38650 207590 38850
rect 207910 38650 207980 38850
rect 204150 38520 204350 38590
rect 204650 38520 204850 38590
rect 205150 38520 205350 38590
rect 205650 38520 205850 38590
rect 206150 38520 206350 38590
rect 206650 38520 206850 38590
rect 207150 38520 207350 38590
rect 207650 38520 207850 38590
rect 204150 38410 204350 38480
rect 204650 38410 204850 38480
rect 205150 38410 205350 38480
rect 205650 38410 205850 38480
rect 206150 38410 206350 38480
rect 206650 38410 206850 38480
rect 207150 38410 207350 38480
rect 207650 38410 207850 38480
rect 204020 38150 204090 38350
rect 204410 38150 204480 38350
rect 204520 38150 204590 38350
rect 204910 38150 204980 38350
rect 205020 38150 205090 38350
rect 205410 38150 205480 38350
rect 205520 38150 205590 38350
rect 205910 38150 205980 38350
rect 206020 38150 206090 38350
rect 206410 38150 206480 38350
rect 206520 38150 206590 38350
rect 206910 38150 206980 38350
rect 207020 38150 207090 38350
rect 207410 38150 207480 38350
rect 207520 38150 207590 38350
rect 207910 38150 207980 38350
rect 204150 38020 204350 38090
rect 204650 38020 204850 38090
rect 205150 38020 205350 38090
rect 205650 38020 205850 38090
rect 206150 38020 206350 38090
rect 206650 38020 206850 38090
rect 207150 38020 207350 38090
rect 207650 38020 207850 38090
rect 204150 37910 204350 37980
rect 204650 37910 204850 37980
rect 205150 37910 205350 37980
rect 205650 37910 205850 37980
rect 206150 37910 206350 37980
rect 206650 37910 206850 37980
rect 207150 37910 207350 37980
rect 207650 37910 207850 37980
rect 204020 37650 204090 37850
rect 204410 37650 204480 37850
rect 204520 37650 204590 37850
rect 204910 37650 204980 37850
rect 205020 37650 205090 37850
rect 205410 37650 205480 37850
rect 205520 37650 205590 37850
rect 205910 37650 205980 37850
rect 206020 37650 206090 37850
rect 206410 37650 206480 37850
rect 206520 37650 206590 37850
rect 206910 37650 206980 37850
rect 207020 37650 207090 37850
rect 207410 37650 207480 37850
rect 207520 37650 207590 37850
rect 207910 37650 207980 37850
rect 204150 37520 204350 37590
rect 204650 37520 204850 37590
rect 205150 37520 205350 37590
rect 205650 37520 205850 37590
rect 206150 37520 206350 37590
rect 206650 37520 206850 37590
rect 207150 37520 207350 37590
rect 207650 37520 207850 37590
rect 204150 37410 204350 37480
rect 204650 37410 204850 37480
rect 205150 37410 205350 37480
rect 205650 37410 205850 37480
rect 206150 37410 206350 37480
rect 206650 37410 206850 37480
rect 207150 37410 207350 37480
rect 207650 37410 207850 37480
rect 204020 37150 204090 37350
rect 204410 37150 204480 37350
rect 204520 37150 204590 37350
rect 204910 37150 204980 37350
rect 205020 37150 205090 37350
rect 205410 37150 205480 37350
rect 205520 37150 205590 37350
rect 205910 37150 205980 37350
rect 206020 37150 206090 37350
rect 206410 37150 206480 37350
rect 206520 37150 206590 37350
rect 206910 37150 206980 37350
rect 207020 37150 207090 37350
rect 207410 37150 207480 37350
rect 207520 37150 207590 37350
rect 207910 37150 207980 37350
rect 204150 37020 204350 37090
rect 204650 37020 204850 37090
rect 205150 37020 205350 37090
rect 205650 37020 205850 37090
rect 206150 37020 206350 37090
rect 206650 37020 206850 37090
rect 207150 37020 207350 37090
rect 207650 37020 207850 37090
rect 204150 36910 204350 36980
rect 204650 36910 204850 36980
rect 205150 36910 205350 36980
rect 205650 36910 205850 36980
rect 206150 36910 206350 36980
rect 206650 36910 206850 36980
rect 207150 36910 207350 36980
rect 207650 36910 207850 36980
rect 204020 36650 204090 36850
rect 204410 36650 204480 36850
rect 204520 36650 204590 36850
rect 204910 36650 204980 36850
rect 205020 36650 205090 36850
rect 205410 36650 205480 36850
rect 205520 36650 205590 36850
rect 205910 36650 205980 36850
rect 206020 36650 206090 36850
rect 206410 36650 206480 36850
rect 206520 36650 206590 36850
rect 206910 36650 206980 36850
rect 207020 36650 207090 36850
rect 207410 36650 207480 36850
rect 207520 36650 207590 36850
rect 207910 36650 207980 36850
rect 204150 36520 204350 36590
rect 204650 36520 204850 36590
rect 205150 36520 205350 36590
rect 205650 36520 205850 36590
rect 206150 36520 206350 36590
rect 206650 36520 206850 36590
rect 207150 36520 207350 36590
rect 207650 36520 207850 36590
rect 204150 36410 204350 36480
rect 204650 36410 204850 36480
rect 205150 36410 205350 36480
rect 205650 36410 205850 36480
rect 206150 36410 206350 36480
rect 206650 36410 206850 36480
rect 207150 36410 207350 36480
rect 207650 36410 207850 36480
rect 204020 36150 204090 36350
rect 204410 36150 204480 36350
rect 204520 36150 204590 36350
rect 204910 36150 204980 36350
rect 205020 36150 205090 36350
rect 205410 36150 205480 36350
rect 205520 36150 205590 36350
rect 205910 36150 205980 36350
rect 206020 36150 206090 36350
rect 206410 36150 206480 36350
rect 206520 36150 206590 36350
rect 206910 36150 206980 36350
rect 207020 36150 207090 36350
rect 207410 36150 207480 36350
rect 207520 36150 207590 36350
rect 207910 36150 207980 36350
rect 204150 36020 204350 36090
rect 204650 36020 204850 36090
rect 205150 36020 205350 36090
rect 205650 36020 205850 36090
rect 206150 36020 206350 36090
rect 206650 36020 206850 36090
rect 207150 36020 207350 36090
rect 207650 36020 207850 36090
rect 204150 35910 204350 35980
rect 204650 35910 204850 35980
rect 205150 35910 205350 35980
rect 205650 35910 205850 35980
rect 206150 35910 206350 35980
rect 206650 35910 206850 35980
rect 207150 35910 207350 35980
rect 207650 35910 207850 35980
rect 204020 35650 204090 35850
rect 204410 35650 204480 35850
rect 204520 35650 204590 35850
rect 204910 35650 204980 35850
rect 205020 35650 205090 35850
rect 205410 35650 205480 35850
rect 205520 35650 205590 35850
rect 205910 35650 205980 35850
rect 206020 35650 206090 35850
rect 206410 35650 206480 35850
rect 206520 35650 206590 35850
rect 206910 35650 206980 35850
rect 207020 35650 207090 35850
rect 207410 35650 207480 35850
rect 207520 35650 207590 35850
rect 207910 35650 207980 35850
rect 204150 35520 204350 35590
rect 204650 35520 204850 35590
rect 205150 35520 205350 35590
rect 205650 35520 205850 35590
rect 206150 35520 206350 35590
rect 206650 35520 206850 35590
rect 207150 35520 207350 35590
rect 207650 35520 207850 35590
rect 204150 35410 204350 35480
rect 204650 35410 204850 35480
rect 205150 35410 205350 35480
rect 205650 35410 205850 35480
rect 206150 35410 206350 35480
rect 206650 35410 206850 35480
rect 207150 35410 207350 35480
rect 207650 35410 207850 35480
rect 204020 35150 204090 35350
rect 204410 35150 204480 35350
rect 204520 35150 204590 35350
rect 204910 35150 204980 35350
rect 205020 35150 205090 35350
rect 205410 35150 205480 35350
rect 205520 35150 205590 35350
rect 205910 35150 205980 35350
rect 206020 35150 206090 35350
rect 206410 35150 206480 35350
rect 206520 35150 206590 35350
rect 206910 35150 206980 35350
rect 207020 35150 207090 35350
rect 207410 35150 207480 35350
rect 207520 35150 207590 35350
rect 207910 35150 207980 35350
rect 204150 35020 204350 35090
rect 204650 35020 204850 35090
rect 205150 35020 205350 35090
rect 205650 35020 205850 35090
rect 206150 35020 206350 35090
rect 206650 35020 206850 35090
rect 207150 35020 207350 35090
rect 207650 35020 207850 35090
rect 204150 34910 204350 34980
rect 204650 34910 204850 34980
rect 205150 34910 205350 34980
rect 205650 34910 205850 34980
rect 206150 34910 206350 34980
rect 206650 34910 206850 34980
rect 207150 34910 207350 34980
rect 207650 34910 207850 34980
rect 204020 34650 204090 34850
rect 204410 34650 204480 34850
rect 204520 34650 204590 34850
rect 204910 34650 204980 34850
rect 205020 34650 205090 34850
rect 205410 34650 205480 34850
rect 205520 34650 205590 34850
rect 205910 34650 205980 34850
rect 206020 34650 206090 34850
rect 206410 34650 206480 34850
rect 206520 34650 206590 34850
rect 206910 34650 206980 34850
rect 207020 34650 207090 34850
rect 207410 34650 207480 34850
rect 207520 34650 207590 34850
rect 207910 34650 207980 34850
rect 204150 34520 204350 34590
rect 204650 34520 204850 34590
rect 205150 34520 205350 34590
rect 205650 34520 205850 34590
rect 206150 34520 206350 34590
rect 206650 34520 206850 34590
rect 207150 34520 207350 34590
rect 207650 34520 207850 34590
rect 204150 34410 204350 34480
rect 204650 34410 204850 34480
rect 205150 34410 205350 34480
rect 205650 34410 205850 34480
rect 206150 34410 206350 34480
rect 206650 34410 206850 34480
rect 207150 34410 207350 34480
rect 207650 34410 207850 34480
rect 204020 34150 204090 34350
rect 204410 34150 204480 34350
rect 204520 34150 204590 34350
rect 204910 34150 204980 34350
rect 205020 34150 205090 34350
rect 205410 34150 205480 34350
rect 205520 34150 205590 34350
rect 205910 34150 205980 34350
rect 206020 34150 206090 34350
rect 206410 34150 206480 34350
rect 206520 34150 206590 34350
rect 206910 34150 206980 34350
rect 207020 34150 207090 34350
rect 207410 34150 207480 34350
rect 207520 34150 207590 34350
rect 207910 34150 207980 34350
rect 204150 34020 204350 34090
rect 204650 34020 204850 34090
rect 205150 34020 205350 34090
rect 205650 34020 205850 34090
rect 206150 34020 206350 34090
rect 206650 34020 206850 34090
rect 207150 34020 207350 34090
rect 207650 34020 207850 34090
rect 204150 33910 204350 33980
rect 204650 33910 204850 33980
rect 205150 33910 205350 33980
rect 205650 33910 205850 33980
rect 206150 33910 206350 33980
rect 206650 33910 206850 33980
rect 207150 33910 207350 33980
rect 207650 33910 207850 33980
rect 204020 33650 204090 33850
rect 204410 33650 204480 33850
rect 204520 33650 204590 33850
rect 204910 33650 204980 33850
rect 205020 33650 205090 33850
rect 205410 33650 205480 33850
rect 205520 33650 205590 33850
rect 205910 33650 205980 33850
rect 206020 33650 206090 33850
rect 206410 33650 206480 33850
rect 206520 33650 206590 33850
rect 206910 33650 206980 33850
rect 207020 33650 207090 33850
rect 207410 33650 207480 33850
rect 207520 33650 207590 33850
rect 207910 33650 207980 33850
rect 204150 33520 204350 33590
rect 204650 33520 204850 33590
rect 205150 33520 205350 33590
rect 205650 33520 205850 33590
rect 206150 33520 206350 33590
rect 206650 33520 206850 33590
rect 207150 33520 207350 33590
rect 207650 33520 207850 33590
rect 204150 33410 204350 33480
rect 204650 33410 204850 33480
rect 205150 33410 205350 33480
rect 205650 33410 205850 33480
rect 206150 33410 206350 33480
rect 206650 33410 206850 33480
rect 207150 33410 207350 33480
rect 207650 33410 207850 33480
rect 204020 33150 204090 33350
rect 204410 33150 204480 33350
rect 204520 33150 204590 33350
rect 204910 33150 204980 33350
rect 205020 33150 205090 33350
rect 205410 33150 205480 33350
rect 205520 33150 205590 33350
rect 205910 33150 205980 33350
rect 206020 33150 206090 33350
rect 206410 33150 206480 33350
rect 206520 33150 206590 33350
rect 206910 33150 206980 33350
rect 207020 33150 207090 33350
rect 207410 33150 207480 33350
rect 207520 33150 207590 33350
rect 207910 33150 207980 33350
rect 204150 33020 204350 33090
rect 204650 33020 204850 33090
rect 205150 33020 205350 33090
rect 205650 33020 205850 33090
rect 206150 33020 206350 33090
rect 206650 33020 206850 33090
rect 207150 33020 207350 33090
rect 207650 33020 207850 33090
rect 204150 32910 204350 32980
rect 204650 32910 204850 32980
rect 205150 32910 205350 32980
rect 205650 32910 205850 32980
rect 206150 32910 206350 32980
rect 206650 32910 206850 32980
rect 207150 32910 207350 32980
rect 207650 32910 207850 32980
rect 204020 32650 204090 32850
rect 204410 32650 204480 32850
rect 204520 32650 204590 32850
rect 204910 32650 204980 32850
rect 205020 32650 205090 32850
rect 205410 32650 205480 32850
rect 205520 32650 205590 32850
rect 205910 32650 205980 32850
rect 206020 32650 206090 32850
rect 206410 32650 206480 32850
rect 206520 32650 206590 32850
rect 206910 32650 206980 32850
rect 207020 32650 207090 32850
rect 207410 32650 207480 32850
rect 207520 32650 207590 32850
rect 207910 32650 207980 32850
rect 204150 32520 204350 32590
rect 204650 32520 204850 32590
rect 205150 32520 205350 32590
rect 205650 32520 205850 32590
rect 206150 32520 206350 32590
rect 206650 32520 206850 32590
rect 207150 32520 207350 32590
rect 207650 32520 207850 32590
rect 204150 32410 204350 32480
rect 204650 32410 204850 32480
rect 205150 32410 205350 32480
rect 205650 32410 205850 32480
rect 206150 32410 206350 32480
rect 206650 32410 206850 32480
rect 207150 32410 207350 32480
rect 207650 32410 207850 32480
rect 204020 32150 204090 32350
rect 204410 32150 204480 32350
rect 204520 32150 204590 32350
rect 204910 32150 204980 32350
rect 205020 32150 205090 32350
rect 205410 32150 205480 32350
rect 205520 32150 205590 32350
rect 205910 32150 205980 32350
rect 206020 32150 206090 32350
rect 206410 32150 206480 32350
rect 206520 32150 206590 32350
rect 206910 32150 206980 32350
rect 207020 32150 207090 32350
rect 207410 32150 207480 32350
rect 207520 32150 207590 32350
rect 207910 32150 207980 32350
rect 204150 32020 204350 32090
rect 204650 32020 204850 32090
rect 205150 32020 205350 32090
rect 205650 32020 205850 32090
rect 206150 32020 206350 32090
rect 206650 32020 206850 32090
rect 207150 32020 207350 32090
rect 207650 32020 207850 32090
rect 204150 31910 204350 31980
rect 204650 31910 204850 31980
rect 205150 31910 205350 31980
rect 205650 31910 205850 31980
rect 206150 31910 206350 31980
rect 206650 31910 206850 31980
rect 207150 31910 207350 31980
rect 207650 31910 207850 31980
rect 204020 31650 204090 31850
rect 204410 31650 204480 31850
rect 204520 31650 204590 31850
rect 204910 31650 204980 31850
rect 205020 31650 205090 31850
rect 205410 31650 205480 31850
rect 205520 31650 205590 31850
rect 205910 31650 205980 31850
rect 206020 31650 206090 31850
rect 206410 31650 206480 31850
rect 206520 31650 206590 31850
rect 206910 31650 206980 31850
rect 207020 31650 207090 31850
rect 207410 31650 207480 31850
rect 207520 31650 207590 31850
rect 207910 31650 207980 31850
rect 204150 31520 204350 31590
rect 204650 31520 204850 31590
rect 205150 31520 205350 31590
rect 205650 31520 205850 31590
rect 206150 31520 206350 31590
rect 206650 31520 206850 31590
rect 207150 31520 207350 31590
rect 207650 31520 207850 31590
rect 204150 31410 204350 31480
rect 204650 31410 204850 31480
rect 205150 31410 205350 31480
rect 205650 31410 205850 31480
rect 206150 31410 206350 31480
rect 206650 31410 206850 31480
rect 207150 31410 207350 31480
rect 207650 31410 207850 31480
rect 204020 31150 204090 31350
rect 204410 31150 204480 31350
rect 204520 31150 204590 31350
rect 204910 31150 204980 31350
rect 205020 31150 205090 31350
rect 205410 31150 205480 31350
rect 205520 31150 205590 31350
rect 205910 31150 205980 31350
rect 206020 31150 206090 31350
rect 206410 31150 206480 31350
rect 206520 31150 206590 31350
rect 206910 31150 206980 31350
rect 207020 31150 207090 31350
rect 207410 31150 207480 31350
rect 207520 31150 207590 31350
rect 207910 31150 207980 31350
rect 204150 31020 204350 31090
rect 204650 31020 204850 31090
rect 205150 31020 205350 31090
rect 205650 31020 205850 31090
rect 206150 31020 206350 31090
rect 206650 31020 206850 31090
rect 207150 31020 207350 31090
rect 207650 31020 207850 31090
rect 204150 30910 204350 30980
rect 204650 30910 204850 30980
rect 205150 30910 205350 30980
rect 205650 30910 205850 30980
rect 206150 30910 206350 30980
rect 206650 30910 206850 30980
rect 207150 30910 207350 30980
rect 207650 30910 207850 30980
rect 204020 30650 204090 30850
rect 204410 30650 204480 30850
rect 204520 30650 204590 30850
rect 204910 30650 204980 30850
rect 205020 30650 205090 30850
rect 205410 30650 205480 30850
rect 205520 30650 205590 30850
rect 205910 30650 205980 30850
rect 206020 30650 206090 30850
rect 206410 30650 206480 30850
rect 206520 30650 206590 30850
rect 206910 30650 206980 30850
rect 207020 30650 207090 30850
rect 207410 30650 207480 30850
rect 207520 30650 207590 30850
rect 207910 30650 207980 30850
rect 204150 30520 204350 30590
rect 204650 30520 204850 30590
rect 205150 30520 205350 30590
rect 205650 30520 205850 30590
rect 206150 30520 206350 30590
rect 206650 30520 206850 30590
rect 207150 30520 207350 30590
rect 207650 30520 207850 30590
rect 204150 30410 204350 30480
rect 204650 30410 204850 30480
rect 205150 30410 205350 30480
rect 205650 30410 205850 30480
rect 206150 30410 206350 30480
rect 206650 30410 206850 30480
rect 207150 30410 207350 30480
rect 207650 30410 207850 30480
rect 204020 30150 204090 30350
rect 204410 30150 204480 30350
rect 204520 30150 204590 30350
rect 204910 30150 204980 30350
rect 205020 30150 205090 30350
rect 205410 30150 205480 30350
rect 205520 30150 205590 30350
rect 205910 30150 205980 30350
rect 206020 30150 206090 30350
rect 206410 30150 206480 30350
rect 206520 30150 206590 30350
rect 206910 30150 206980 30350
rect 207020 30150 207090 30350
rect 207410 30150 207480 30350
rect 207520 30150 207590 30350
rect 207910 30150 207980 30350
rect 204150 30020 204350 30090
rect 204650 30020 204850 30090
rect 205150 30020 205350 30090
rect 205650 30020 205850 30090
rect 206150 30020 206350 30090
rect 206650 30020 206850 30090
rect 207150 30020 207350 30090
rect 207650 30020 207850 30090
rect 204150 29910 204350 29980
rect 204650 29910 204850 29980
rect 205150 29910 205350 29980
rect 205650 29910 205850 29980
rect 206150 29910 206350 29980
rect 206650 29910 206850 29980
rect 207150 29910 207350 29980
rect 207650 29910 207850 29980
rect 204020 29650 204090 29850
rect 204410 29650 204480 29850
rect 204520 29650 204590 29850
rect 204910 29650 204980 29850
rect 205020 29650 205090 29850
rect 205410 29650 205480 29850
rect 205520 29650 205590 29850
rect 205910 29650 205980 29850
rect 206020 29650 206090 29850
rect 206410 29650 206480 29850
rect 206520 29650 206590 29850
rect 206910 29650 206980 29850
rect 207020 29650 207090 29850
rect 207410 29650 207480 29850
rect 207520 29650 207590 29850
rect 207910 29650 207980 29850
rect 204150 29520 204350 29590
rect 204650 29520 204850 29590
rect 205150 29520 205350 29590
rect 205650 29520 205850 29590
rect 206150 29520 206350 29590
rect 206650 29520 206850 29590
rect 207150 29520 207350 29590
rect 207650 29520 207850 29590
rect 204150 29410 204350 29480
rect 204650 29410 204850 29480
rect 205150 29410 205350 29480
rect 205650 29410 205850 29480
rect 206150 29410 206350 29480
rect 206650 29410 206850 29480
rect 207150 29410 207350 29480
rect 207650 29410 207850 29480
rect 204020 29150 204090 29350
rect 204410 29150 204480 29350
rect 204520 29150 204590 29350
rect 204910 29150 204980 29350
rect 205020 29150 205090 29350
rect 205410 29150 205480 29350
rect 205520 29150 205590 29350
rect 205910 29150 205980 29350
rect 206020 29150 206090 29350
rect 206410 29150 206480 29350
rect 206520 29150 206590 29350
rect 206910 29150 206980 29350
rect 207020 29150 207090 29350
rect 207410 29150 207480 29350
rect 207520 29150 207590 29350
rect 207910 29150 207980 29350
rect 204150 29020 204350 29090
rect 204650 29020 204850 29090
rect 205150 29020 205350 29090
rect 205650 29020 205850 29090
rect 206150 29020 206350 29090
rect 206650 29020 206850 29090
rect 207150 29020 207350 29090
rect 207650 29020 207850 29090
rect 204150 28910 204350 28980
rect 204650 28910 204850 28980
rect 205150 28910 205350 28980
rect 205650 28910 205850 28980
rect 206150 28910 206350 28980
rect 206650 28910 206850 28980
rect 207150 28910 207350 28980
rect 207650 28910 207850 28980
rect 204020 28650 204090 28850
rect 204410 28650 204480 28850
rect 204520 28650 204590 28850
rect 204910 28650 204980 28850
rect 205020 28650 205090 28850
rect 205410 28650 205480 28850
rect 205520 28650 205590 28850
rect 205910 28650 205980 28850
rect 206020 28650 206090 28850
rect 206410 28650 206480 28850
rect 206520 28650 206590 28850
rect 206910 28650 206980 28850
rect 207020 28650 207090 28850
rect 207410 28650 207480 28850
rect 207520 28650 207590 28850
rect 207910 28650 207980 28850
rect 204150 28520 204350 28590
rect 204650 28520 204850 28590
rect 205150 28520 205350 28590
rect 205650 28520 205850 28590
rect 206150 28520 206350 28590
rect 206650 28520 206850 28590
rect 207150 28520 207350 28590
rect 207650 28520 207850 28590
rect 204150 28410 204350 28480
rect 204650 28410 204850 28480
rect 205150 28410 205350 28480
rect 205650 28410 205850 28480
rect 206150 28410 206350 28480
rect 206650 28410 206850 28480
rect 207150 28410 207350 28480
rect 207650 28410 207850 28480
rect 204020 28150 204090 28350
rect 204410 28150 204480 28350
rect 204520 28150 204590 28350
rect 204910 28150 204980 28350
rect 205020 28150 205090 28350
rect 205410 28150 205480 28350
rect 205520 28150 205590 28350
rect 205910 28150 205980 28350
rect 206020 28150 206090 28350
rect 206410 28150 206480 28350
rect 206520 28150 206590 28350
rect 206910 28150 206980 28350
rect 207020 28150 207090 28350
rect 207410 28150 207480 28350
rect 207520 28150 207590 28350
rect 207910 28150 207980 28350
rect 204150 28020 204350 28090
rect 204650 28020 204850 28090
rect 205150 28020 205350 28090
rect 205650 28020 205850 28090
rect 206150 28020 206350 28090
rect 206650 28020 206850 28090
rect 207150 28020 207350 28090
rect 207650 28020 207850 28090
rect 204150 27910 204350 27980
rect 204650 27910 204850 27980
rect 205150 27910 205350 27980
rect 205650 27910 205850 27980
rect 206150 27910 206350 27980
rect 206650 27910 206850 27980
rect 207150 27910 207350 27980
rect 207650 27910 207850 27980
rect 204020 27650 204090 27850
rect 204410 27650 204480 27850
rect 204520 27650 204590 27850
rect 204910 27650 204980 27850
rect 205020 27650 205090 27850
rect 205410 27650 205480 27850
rect 205520 27650 205590 27850
rect 205910 27650 205980 27850
rect 206020 27650 206090 27850
rect 206410 27650 206480 27850
rect 206520 27650 206590 27850
rect 206910 27650 206980 27850
rect 207020 27650 207090 27850
rect 207410 27650 207480 27850
rect 207520 27650 207590 27850
rect 207910 27650 207980 27850
rect 204150 27520 204350 27590
rect 204650 27520 204850 27590
rect 205150 27520 205350 27590
rect 205650 27520 205850 27590
rect 206150 27520 206350 27590
rect 206650 27520 206850 27590
rect 207150 27520 207350 27590
rect 207650 27520 207850 27590
rect 204150 27410 204350 27480
rect 204650 27410 204850 27480
rect 205150 27410 205350 27480
rect 205650 27410 205850 27480
rect 206150 27410 206350 27480
rect 206650 27410 206850 27480
rect 207150 27410 207350 27480
rect 207650 27410 207850 27480
rect 204020 27150 204090 27350
rect 204410 27150 204480 27350
rect 204520 27150 204590 27350
rect 204910 27150 204980 27350
rect 205020 27150 205090 27350
rect 205410 27150 205480 27350
rect 205520 27150 205590 27350
rect 205910 27150 205980 27350
rect 206020 27150 206090 27350
rect 206410 27150 206480 27350
rect 206520 27150 206590 27350
rect 206910 27150 206980 27350
rect 207020 27150 207090 27350
rect 207410 27150 207480 27350
rect 207520 27150 207590 27350
rect 207910 27150 207980 27350
rect 204150 27020 204350 27090
rect 204650 27020 204850 27090
rect 205150 27020 205350 27090
rect 205650 27020 205850 27090
rect 206150 27020 206350 27090
rect 206650 27020 206850 27090
rect 207150 27020 207350 27090
rect 207650 27020 207850 27090
rect 204150 26910 204350 26980
rect 204650 26910 204850 26980
rect 205150 26910 205350 26980
rect 205650 26910 205850 26980
rect 206150 26910 206350 26980
rect 206650 26910 206850 26980
rect 207150 26910 207350 26980
rect 207650 26910 207850 26980
rect 204020 26650 204090 26850
rect 204410 26650 204480 26850
rect 204520 26650 204590 26850
rect 204910 26650 204980 26850
rect 205020 26650 205090 26850
rect 205410 26650 205480 26850
rect 205520 26650 205590 26850
rect 205910 26650 205980 26850
rect 206020 26650 206090 26850
rect 206410 26650 206480 26850
rect 206520 26650 206590 26850
rect 206910 26650 206980 26850
rect 207020 26650 207090 26850
rect 207410 26650 207480 26850
rect 207520 26650 207590 26850
rect 207910 26650 207980 26850
rect 204150 26520 204350 26590
rect 204650 26520 204850 26590
rect 205150 26520 205350 26590
rect 205650 26520 205850 26590
rect 206150 26520 206350 26590
rect 206650 26520 206850 26590
rect 207150 26520 207350 26590
rect 207650 26520 207850 26590
rect 204150 26410 204350 26480
rect 204650 26410 204850 26480
rect 205150 26410 205350 26480
rect 205650 26410 205850 26480
rect 206150 26410 206350 26480
rect 206650 26410 206850 26480
rect 207150 26410 207350 26480
rect 207650 26410 207850 26480
rect 204020 26150 204090 26350
rect 204410 26150 204480 26350
rect 204520 26150 204590 26350
rect 204910 26150 204980 26350
rect 205020 26150 205090 26350
rect 205410 26150 205480 26350
rect 205520 26150 205590 26350
rect 205910 26150 205980 26350
rect 206020 26150 206090 26350
rect 206410 26150 206480 26350
rect 206520 26150 206590 26350
rect 206910 26150 206980 26350
rect 207020 26150 207090 26350
rect 207410 26150 207480 26350
rect 207520 26150 207590 26350
rect 207910 26150 207980 26350
rect 204150 26020 204350 26090
rect 204650 26020 204850 26090
rect 205150 26020 205350 26090
rect 205650 26020 205850 26090
rect 206150 26020 206350 26090
rect 206650 26020 206850 26090
rect 207150 26020 207350 26090
rect 207650 26020 207850 26090
rect 204150 25910 204350 25980
rect 204650 25910 204850 25980
rect 205150 25910 205350 25980
rect 205650 25910 205850 25980
rect 206150 25910 206350 25980
rect 206650 25910 206850 25980
rect 207150 25910 207350 25980
rect 207650 25910 207850 25980
rect 204020 25650 204090 25850
rect 204410 25650 204480 25850
rect 204520 25650 204590 25850
rect 204910 25650 204980 25850
rect 205020 25650 205090 25850
rect 205410 25650 205480 25850
rect 205520 25650 205590 25850
rect 205910 25650 205980 25850
rect 206020 25650 206090 25850
rect 206410 25650 206480 25850
rect 206520 25650 206590 25850
rect 206910 25650 206980 25850
rect 207020 25650 207090 25850
rect 207410 25650 207480 25850
rect 207520 25650 207590 25850
rect 207910 25650 207980 25850
rect 204150 25520 204350 25590
rect 204650 25520 204850 25590
rect 205150 25520 205350 25590
rect 205650 25520 205850 25590
rect 206150 25520 206350 25590
rect 206650 25520 206850 25590
rect 207150 25520 207350 25590
rect 207650 25520 207850 25590
rect 204150 25410 204350 25480
rect 204650 25410 204850 25480
rect 205150 25410 205350 25480
rect 205650 25410 205850 25480
rect 206150 25410 206350 25480
rect 206650 25410 206850 25480
rect 207150 25410 207350 25480
rect 207650 25410 207850 25480
rect 204020 25150 204090 25350
rect 204410 25150 204480 25350
rect 204520 25150 204590 25350
rect 204910 25150 204980 25350
rect 205020 25150 205090 25350
rect 205410 25150 205480 25350
rect 205520 25150 205590 25350
rect 205910 25150 205980 25350
rect 206020 25150 206090 25350
rect 206410 25150 206480 25350
rect 206520 25150 206590 25350
rect 206910 25150 206980 25350
rect 207020 25150 207090 25350
rect 207410 25150 207480 25350
rect 207520 25150 207590 25350
rect 207910 25150 207980 25350
rect 204150 25020 204350 25090
rect 204650 25020 204850 25090
rect 205150 25020 205350 25090
rect 205650 25020 205850 25090
rect 206150 25020 206350 25090
rect 206650 25020 206850 25090
rect 207150 25020 207350 25090
rect 207650 25020 207850 25090
rect 204150 24910 204350 24980
rect 204650 24910 204850 24980
rect 205150 24910 205350 24980
rect 205650 24910 205850 24980
rect 206150 24910 206350 24980
rect 206650 24910 206850 24980
rect 207150 24910 207350 24980
rect 207650 24910 207850 24980
rect 204020 24650 204090 24850
rect 204410 24650 204480 24850
rect 204520 24650 204590 24850
rect 204910 24650 204980 24850
rect 205020 24650 205090 24850
rect 205410 24650 205480 24850
rect 205520 24650 205590 24850
rect 205910 24650 205980 24850
rect 206020 24650 206090 24850
rect 206410 24650 206480 24850
rect 206520 24650 206590 24850
rect 206910 24650 206980 24850
rect 207020 24650 207090 24850
rect 207410 24650 207480 24850
rect 207520 24650 207590 24850
rect 207910 24650 207980 24850
rect 204150 24520 204350 24590
rect 204650 24520 204850 24590
rect 205150 24520 205350 24590
rect 205650 24520 205850 24590
rect 206150 24520 206350 24590
rect 206650 24520 206850 24590
rect 207150 24520 207350 24590
rect 207650 24520 207850 24590
rect 204150 24410 204350 24480
rect 204650 24410 204850 24480
rect 205150 24410 205350 24480
rect 205650 24410 205850 24480
rect 206150 24410 206350 24480
rect 206650 24410 206850 24480
rect 207150 24410 207350 24480
rect 207650 24410 207850 24480
rect 204020 24150 204090 24350
rect 204410 24150 204480 24350
rect 204520 24150 204590 24350
rect 204910 24150 204980 24350
rect 205020 24150 205090 24350
rect 205410 24150 205480 24350
rect 205520 24150 205590 24350
rect 205910 24150 205980 24350
rect 206020 24150 206090 24350
rect 206410 24150 206480 24350
rect 206520 24150 206590 24350
rect 206910 24150 206980 24350
rect 207020 24150 207090 24350
rect 207410 24150 207480 24350
rect 207520 24150 207590 24350
rect 207910 24150 207980 24350
rect 204150 24020 204350 24090
rect 204650 24020 204850 24090
rect 205150 24020 205350 24090
rect 205650 24020 205850 24090
rect 206150 24020 206350 24090
rect 206650 24020 206850 24090
rect 207150 24020 207350 24090
rect 207650 24020 207850 24090
rect 204150 23910 204350 23980
rect 204650 23910 204850 23980
rect 205150 23910 205350 23980
rect 205650 23910 205850 23980
rect 206150 23910 206350 23980
rect 206650 23910 206850 23980
rect 207150 23910 207350 23980
rect 207650 23910 207850 23980
rect 204020 23650 204090 23850
rect 204410 23650 204480 23850
rect 204520 23650 204590 23850
rect 204910 23650 204980 23850
rect 205020 23650 205090 23850
rect 205410 23650 205480 23850
rect 205520 23650 205590 23850
rect 205910 23650 205980 23850
rect 206020 23650 206090 23850
rect 206410 23650 206480 23850
rect 206520 23650 206590 23850
rect 206910 23650 206980 23850
rect 207020 23650 207090 23850
rect 207410 23650 207480 23850
rect 207520 23650 207590 23850
rect 207910 23650 207980 23850
rect 204150 23520 204350 23590
rect 204650 23520 204850 23590
rect 205150 23520 205350 23590
rect 205650 23520 205850 23590
rect 206150 23520 206350 23590
rect 206650 23520 206850 23590
rect 207150 23520 207350 23590
rect 207650 23520 207850 23590
rect 204150 23410 204350 23480
rect 204650 23410 204850 23480
rect 205150 23410 205350 23480
rect 205650 23410 205850 23480
rect 206150 23410 206350 23480
rect 206650 23410 206850 23480
rect 207150 23410 207350 23480
rect 207650 23410 207850 23480
rect 204020 23150 204090 23350
rect 204410 23150 204480 23350
rect 204520 23150 204590 23350
rect 204910 23150 204980 23350
rect 205020 23150 205090 23350
rect 205410 23150 205480 23350
rect 205520 23150 205590 23350
rect 205910 23150 205980 23350
rect 206020 23150 206090 23350
rect 206410 23150 206480 23350
rect 206520 23150 206590 23350
rect 206910 23150 206980 23350
rect 207020 23150 207090 23350
rect 207410 23150 207480 23350
rect 207520 23150 207590 23350
rect 207910 23150 207980 23350
rect 204150 23020 204350 23090
rect 204650 23020 204850 23090
rect 205150 23020 205350 23090
rect 205650 23020 205850 23090
rect 206150 23020 206350 23090
rect 206650 23020 206850 23090
rect 207150 23020 207350 23090
rect 207650 23020 207850 23090
rect 204150 22910 204350 22980
rect 204650 22910 204850 22980
rect 205150 22910 205350 22980
rect 205650 22910 205850 22980
rect 206150 22910 206350 22980
rect 206650 22910 206850 22980
rect 207150 22910 207350 22980
rect 207650 22910 207850 22980
rect 204020 22650 204090 22850
rect 204410 22650 204480 22850
rect 204520 22650 204590 22850
rect 204910 22650 204980 22850
rect 205020 22650 205090 22850
rect 205410 22650 205480 22850
rect 205520 22650 205590 22850
rect 205910 22650 205980 22850
rect 206020 22650 206090 22850
rect 206410 22650 206480 22850
rect 206520 22650 206590 22850
rect 206910 22650 206980 22850
rect 207020 22650 207090 22850
rect 207410 22650 207480 22850
rect 207520 22650 207590 22850
rect 207910 22650 207980 22850
rect 204150 22520 204350 22590
rect 204650 22520 204850 22590
rect 205150 22520 205350 22590
rect 205650 22520 205850 22590
rect 206150 22520 206350 22590
rect 206650 22520 206850 22590
rect 207150 22520 207350 22590
rect 207650 22520 207850 22590
rect 204150 22410 204350 22480
rect 204650 22410 204850 22480
rect 205150 22410 205350 22480
rect 205650 22410 205850 22480
rect 206150 22410 206350 22480
rect 206650 22410 206850 22480
rect 207150 22410 207350 22480
rect 207650 22410 207850 22480
rect 204020 22150 204090 22350
rect 204410 22150 204480 22350
rect 204520 22150 204590 22350
rect 204910 22150 204980 22350
rect 205020 22150 205090 22350
rect 205410 22150 205480 22350
rect 205520 22150 205590 22350
rect 205910 22150 205980 22350
rect 206020 22150 206090 22350
rect 206410 22150 206480 22350
rect 206520 22150 206590 22350
rect 206910 22150 206980 22350
rect 207020 22150 207090 22350
rect 207410 22150 207480 22350
rect 207520 22150 207590 22350
rect 207910 22150 207980 22350
rect 204150 22020 204350 22090
rect 204650 22020 204850 22090
rect 205150 22020 205350 22090
rect 205650 22020 205850 22090
rect 206150 22020 206350 22090
rect 206650 22020 206850 22090
rect 207150 22020 207350 22090
rect 207650 22020 207850 22090
rect 204150 21910 204350 21980
rect 204650 21910 204850 21980
rect 205150 21910 205350 21980
rect 205650 21910 205850 21980
rect 206150 21910 206350 21980
rect 206650 21910 206850 21980
rect 207150 21910 207350 21980
rect 207650 21910 207850 21980
rect 204020 21650 204090 21850
rect 204410 21650 204480 21850
rect 204520 21650 204590 21850
rect 204910 21650 204980 21850
rect 205020 21650 205090 21850
rect 205410 21650 205480 21850
rect 205520 21650 205590 21850
rect 205910 21650 205980 21850
rect 206020 21650 206090 21850
rect 206410 21650 206480 21850
rect 206520 21650 206590 21850
rect 206910 21650 206980 21850
rect 207020 21650 207090 21850
rect 207410 21650 207480 21850
rect 207520 21650 207590 21850
rect 207910 21650 207980 21850
rect 204150 21520 204350 21590
rect 204650 21520 204850 21590
rect 205150 21520 205350 21590
rect 205650 21520 205850 21590
rect 206150 21520 206350 21590
rect 206650 21520 206850 21590
rect 207150 21520 207350 21590
rect 207650 21520 207850 21590
rect 204150 21410 204350 21480
rect 204650 21410 204850 21480
rect 205150 21410 205350 21480
rect 205650 21410 205850 21480
rect 206150 21410 206350 21480
rect 206650 21410 206850 21480
rect 207150 21410 207350 21480
rect 207650 21410 207850 21480
rect 204020 21150 204090 21350
rect 204410 21150 204480 21350
rect 204520 21150 204590 21350
rect 204910 21150 204980 21350
rect 205020 21150 205090 21350
rect 205410 21150 205480 21350
rect 205520 21150 205590 21350
rect 205910 21150 205980 21350
rect 206020 21150 206090 21350
rect 206410 21150 206480 21350
rect 206520 21150 206590 21350
rect 206910 21150 206980 21350
rect 207020 21150 207090 21350
rect 207410 21150 207480 21350
rect 207520 21150 207590 21350
rect 207910 21150 207980 21350
rect 204150 21020 204350 21090
rect 204650 21020 204850 21090
rect 205150 21020 205350 21090
rect 205650 21020 205850 21090
rect 206150 21020 206350 21090
rect 206650 21020 206850 21090
rect 207150 21020 207350 21090
rect 207650 21020 207850 21090
rect 204150 20910 204350 20980
rect 204650 20910 204850 20980
rect 205150 20910 205350 20980
rect 205650 20910 205850 20980
rect 206150 20910 206350 20980
rect 206650 20910 206850 20980
rect 207150 20910 207350 20980
rect 207650 20910 207850 20980
rect 204020 20650 204090 20850
rect 204410 20650 204480 20850
rect 204520 20650 204590 20850
rect 204910 20650 204980 20850
rect 205020 20650 205090 20850
rect 205410 20650 205480 20850
rect 205520 20650 205590 20850
rect 205910 20650 205980 20850
rect 206020 20650 206090 20850
rect 206410 20650 206480 20850
rect 206520 20650 206590 20850
rect 206910 20650 206980 20850
rect 207020 20650 207090 20850
rect 207410 20650 207480 20850
rect 207520 20650 207590 20850
rect 207910 20650 207980 20850
rect 204150 20520 204350 20590
rect 204650 20520 204850 20590
rect 205150 20520 205350 20590
rect 205650 20520 205850 20590
rect 206150 20520 206350 20590
rect 206650 20520 206850 20590
rect 207150 20520 207350 20590
rect 207650 20520 207850 20590
rect 204150 20410 204350 20480
rect 204650 20410 204850 20480
rect 205150 20410 205350 20480
rect 205650 20410 205850 20480
rect 206150 20410 206350 20480
rect 206650 20410 206850 20480
rect 207150 20410 207350 20480
rect 207650 20410 207850 20480
rect 204020 20150 204090 20350
rect 204410 20150 204480 20350
rect 204520 20150 204590 20350
rect 204910 20150 204980 20350
rect 205020 20150 205090 20350
rect 205410 20150 205480 20350
rect 205520 20150 205590 20350
rect 205910 20150 205980 20350
rect 206020 20150 206090 20350
rect 206410 20150 206480 20350
rect 206520 20150 206590 20350
rect 206910 20150 206980 20350
rect 207020 20150 207090 20350
rect 207410 20150 207480 20350
rect 207520 20150 207590 20350
rect 207910 20150 207980 20350
rect 204150 20020 204350 20090
rect 204650 20020 204850 20090
rect 205150 20020 205350 20090
rect 205650 20020 205850 20090
rect 206150 20020 206350 20090
rect 206650 20020 206850 20090
rect 207150 20020 207350 20090
rect 207650 20020 207850 20090
rect 204150 19910 204350 19980
rect 204650 19910 204850 19980
rect 205150 19910 205350 19980
rect 205650 19910 205850 19980
rect 206150 19910 206350 19980
rect 206650 19910 206850 19980
rect 207150 19910 207350 19980
rect 207650 19910 207850 19980
rect 204020 19650 204090 19850
rect 204410 19650 204480 19850
rect 204520 19650 204590 19850
rect 204910 19650 204980 19850
rect 205020 19650 205090 19850
rect 205410 19650 205480 19850
rect 205520 19650 205590 19850
rect 205910 19650 205980 19850
rect 206020 19650 206090 19850
rect 206410 19650 206480 19850
rect 206520 19650 206590 19850
rect 206910 19650 206980 19850
rect 207020 19650 207090 19850
rect 207410 19650 207480 19850
rect 207520 19650 207590 19850
rect 207910 19650 207980 19850
rect 204150 19520 204350 19590
rect 204650 19520 204850 19590
rect 205150 19520 205350 19590
rect 205650 19520 205850 19590
rect 206150 19520 206350 19590
rect 206650 19520 206850 19590
rect 207150 19520 207350 19590
rect 207650 19520 207850 19590
rect 204150 19410 204350 19480
rect 204650 19410 204850 19480
rect 205150 19410 205350 19480
rect 205650 19410 205850 19480
rect 206150 19410 206350 19480
rect 206650 19410 206850 19480
rect 207150 19410 207350 19480
rect 207650 19410 207850 19480
rect 204020 19150 204090 19350
rect 204410 19150 204480 19350
rect 204520 19150 204590 19350
rect 204910 19150 204980 19350
rect 205020 19150 205090 19350
rect 205410 19150 205480 19350
rect 205520 19150 205590 19350
rect 205910 19150 205980 19350
rect 206020 19150 206090 19350
rect 206410 19150 206480 19350
rect 206520 19150 206590 19350
rect 206910 19150 206980 19350
rect 207020 19150 207090 19350
rect 207410 19150 207480 19350
rect 207520 19150 207590 19350
rect 207910 19150 207980 19350
rect 204150 19020 204350 19090
rect 204650 19020 204850 19090
rect 205150 19020 205350 19090
rect 205650 19020 205850 19090
rect 206150 19020 206350 19090
rect 206650 19020 206850 19090
rect 207150 19020 207350 19090
rect 207650 19020 207850 19090
rect 204150 18910 204350 18980
rect 204650 18910 204850 18980
rect 205150 18910 205350 18980
rect 205650 18910 205850 18980
rect 206150 18910 206350 18980
rect 206650 18910 206850 18980
rect 207150 18910 207350 18980
rect 207650 18910 207850 18980
rect 204020 18650 204090 18850
rect 204410 18650 204480 18850
rect 204520 18650 204590 18850
rect 204910 18650 204980 18850
rect 205020 18650 205090 18850
rect 205410 18650 205480 18850
rect 205520 18650 205590 18850
rect 205910 18650 205980 18850
rect 206020 18650 206090 18850
rect 206410 18650 206480 18850
rect 206520 18650 206590 18850
rect 206910 18650 206980 18850
rect 207020 18650 207090 18850
rect 207410 18650 207480 18850
rect 207520 18650 207590 18850
rect 207910 18650 207980 18850
rect 204150 18520 204350 18590
rect 204650 18520 204850 18590
rect 205150 18520 205350 18590
rect 205650 18520 205850 18590
rect 206150 18520 206350 18590
rect 206650 18520 206850 18590
rect 207150 18520 207350 18590
rect 207650 18520 207850 18590
rect 204150 18410 204350 18480
rect 204650 18410 204850 18480
rect 205150 18410 205350 18480
rect 205650 18410 205850 18480
rect 206150 18410 206350 18480
rect 206650 18410 206850 18480
rect 207150 18410 207350 18480
rect 207650 18410 207850 18480
rect 204020 18150 204090 18350
rect 204410 18150 204480 18350
rect 204520 18150 204590 18350
rect 204910 18150 204980 18350
rect 205020 18150 205090 18350
rect 205410 18150 205480 18350
rect 205520 18150 205590 18350
rect 205910 18150 205980 18350
rect 206020 18150 206090 18350
rect 206410 18150 206480 18350
rect 206520 18150 206590 18350
rect 206910 18150 206980 18350
rect 207020 18150 207090 18350
rect 207410 18150 207480 18350
rect 207520 18150 207590 18350
rect 207910 18150 207980 18350
rect 204150 18020 204350 18090
rect 204650 18020 204850 18090
rect 205150 18020 205350 18090
rect 205650 18020 205850 18090
rect 206150 18020 206350 18090
rect 206650 18020 206850 18090
rect 207150 18020 207350 18090
rect 207650 18020 207850 18090
rect 204150 17910 204350 17980
rect 204650 17910 204850 17980
rect 205150 17910 205350 17980
rect 205650 17910 205850 17980
rect 206150 17910 206350 17980
rect 206650 17910 206850 17980
rect 207150 17910 207350 17980
rect 207650 17910 207850 17980
rect 204020 17650 204090 17850
rect 204410 17650 204480 17850
rect 204520 17650 204590 17850
rect 204910 17650 204980 17850
rect 205020 17650 205090 17850
rect 205410 17650 205480 17850
rect 205520 17650 205590 17850
rect 205910 17650 205980 17850
rect 206020 17650 206090 17850
rect 206410 17650 206480 17850
rect 206520 17650 206590 17850
rect 206910 17650 206980 17850
rect 207020 17650 207090 17850
rect 207410 17650 207480 17850
rect 207520 17650 207590 17850
rect 207910 17650 207980 17850
rect 204150 17520 204350 17590
rect 204650 17520 204850 17590
rect 205150 17520 205350 17590
rect 205650 17520 205850 17590
rect 206150 17520 206350 17590
rect 206650 17520 206850 17590
rect 207150 17520 207350 17590
rect 207650 17520 207850 17590
rect 204150 17410 204350 17480
rect 204650 17410 204850 17480
rect 205150 17410 205350 17480
rect 205650 17410 205850 17480
rect 206150 17410 206350 17480
rect 206650 17410 206850 17480
rect 207150 17410 207350 17480
rect 207650 17410 207850 17480
rect 204020 17150 204090 17350
rect 204410 17150 204480 17350
rect 204520 17150 204590 17350
rect 204910 17150 204980 17350
rect 205020 17150 205090 17350
rect 205410 17150 205480 17350
rect 205520 17150 205590 17350
rect 205910 17150 205980 17350
rect 206020 17150 206090 17350
rect 206410 17150 206480 17350
rect 206520 17150 206590 17350
rect 206910 17150 206980 17350
rect 207020 17150 207090 17350
rect 207410 17150 207480 17350
rect 207520 17150 207590 17350
rect 207910 17150 207980 17350
rect 204150 17020 204350 17090
rect 204650 17020 204850 17090
rect 205150 17020 205350 17090
rect 205650 17020 205850 17090
rect 206150 17020 206350 17090
rect 206650 17020 206850 17090
rect 207150 17020 207350 17090
rect 207650 17020 207850 17090
rect 204150 16910 204350 16980
rect 204650 16910 204850 16980
rect 205150 16910 205350 16980
rect 205650 16910 205850 16980
rect 206150 16910 206350 16980
rect 206650 16910 206850 16980
rect 207150 16910 207350 16980
rect 207650 16910 207850 16980
rect 204020 16650 204090 16850
rect 204410 16650 204480 16850
rect 204520 16650 204590 16850
rect 204910 16650 204980 16850
rect 205020 16650 205090 16850
rect 205410 16650 205480 16850
rect 205520 16650 205590 16850
rect 205910 16650 205980 16850
rect 206020 16650 206090 16850
rect 206410 16650 206480 16850
rect 206520 16650 206590 16850
rect 206910 16650 206980 16850
rect 207020 16650 207090 16850
rect 207410 16650 207480 16850
rect 207520 16650 207590 16850
rect 207910 16650 207980 16850
rect 204150 16520 204350 16590
rect 204650 16520 204850 16590
rect 205150 16520 205350 16590
rect 205650 16520 205850 16590
rect 206150 16520 206350 16590
rect 206650 16520 206850 16590
rect 207150 16520 207350 16590
rect 207650 16520 207850 16590
rect 204150 16410 204350 16480
rect 204650 16410 204850 16480
rect 205150 16410 205350 16480
rect 205650 16410 205850 16480
rect 206150 16410 206350 16480
rect 206650 16410 206850 16480
rect 207150 16410 207350 16480
rect 207650 16410 207850 16480
rect 204020 16150 204090 16350
rect 204410 16150 204480 16350
rect 204520 16150 204590 16350
rect 204910 16150 204980 16350
rect 205020 16150 205090 16350
rect 205410 16150 205480 16350
rect 205520 16150 205590 16350
rect 205910 16150 205980 16350
rect 206020 16150 206090 16350
rect 206410 16150 206480 16350
rect 206520 16150 206590 16350
rect 206910 16150 206980 16350
rect 207020 16150 207090 16350
rect 207410 16150 207480 16350
rect 207520 16150 207590 16350
rect 207910 16150 207980 16350
rect 204150 16020 204350 16090
rect 204650 16020 204850 16090
rect 205150 16020 205350 16090
rect 205650 16020 205850 16090
rect 206150 16020 206350 16090
rect 206650 16020 206850 16090
rect 207150 16020 207350 16090
rect 207650 16020 207850 16090
rect 204150 15910 204350 15980
rect 204650 15910 204850 15980
rect 205150 15910 205350 15980
rect 205650 15910 205850 15980
rect 206150 15910 206350 15980
rect 206650 15910 206850 15980
rect 207150 15910 207350 15980
rect 207650 15910 207850 15980
rect 204020 15650 204090 15850
rect 204410 15650 204480 15850
rect 204520 15650 204590 15850
rect 204910 15650 204980 15850
rect 205020 15650 205090 15850
rect 205410 15650 205480 15850
rect 205520 15650 205590 15850
rect 205910 15650 205980 15850
rect 206020 15650 206090 15850
rect 206410 15650 206480 15850
rect 206520 15650 206590 15850
rect 206910 15650 206980 15850
rect 207020 15650 207090 15850
rect 207410 15650 207480 15850
rect 207520 15650 207590 15850
rect 207910 15650 207980 15850
rect 204150 15520 204350 15590
rect 204650 15520 204850 15590
rect 205150 15520 205350 15590
rect 205650 15520 205850 15590
rect 206150 15520 206350 15590
rect 206650 15520 206850 15590
rect 207150 15520 207350 15590
rect 207650 15520 207850 15590
rect 204150 15410 204350 15480
rect 204650 15410 204850 15480
rect 205150 15410 205350 15480
rect 205650 15410 205850 15480
rect 206150 15410 206350 15480
rect 206650 15410 206850 15480
rect 207150 15410 207350 15480
rect 207650 15410 207850 15480
rect 204020 15150 204090 15350
rect 204410 15150 204480 15350
rect 204520 15150 204590 15350
rect 204910 15150 204980 15350
rect 205020 15150 205090 15350
rect 205410 15150 205480 15350
rect 205520 15150 205590 15350
rect 205910 15150 205980 15350
rect 206020 15150 206090 15350
rect 206410 15150 206480 15350
rect 206520 15150 206590 15350
rect 206910 15150 206980 15350
rect 207020 15150 207090 15350
rect 207410 15150 207480 15350
rect 207520 15150 207590 15350
rect 207910 15150 207980 15350
rect 204150 15020 204350 15090
rect 204650 15020 204850 15090
rect 205150 15020 205350 15090
rect 205650 15020 205850 15090
rect 206150 15020 206350 15090
rect 206650 15020 206850 15090
rect 207150 15020 207350 15090
rect 207650 15020 207850 15090
rect 204150 14910 204350 14980
rect 204650 14910 204850 14980
rect 205150 14910 205350 14980
rect 205650 14910 205850 14980
rect 206150 14910 206350 14980
rect 206650 14910 206850 14980
rect 207150 14910 207350 14980
rect 207650 14910 207850 14980
rect 204020 14650 204090 14850
rect 204410 14650 204480 14850
rect 204520 14650 204590 14850
rect 204910 14650 204980 14850
rect 205020 14650 205090 14850
rect 205410 14650 205480 14850
rect 205520 14650 205590 14850
rect 205910 14650 205980 14850
rect 206020 14650 206090 14850
rect 206410 14650 206480 14850
rect 206520 14650 206590 14850
rect 206910 14650 206980 14850
rect 207020 14650 207090 14850
rect 207410 14650 207480 14850
rect 207520 14650 207590 14850
rect 207910 14650 207980 14850
rect 204150 14520 204350 14590
rect 204650 14520 204850 14590
rect 205150 14520 205350 14590
rect 205650 14520 205850 14590
rect 206150 14520 206350 14590
rect 206650 14520 206850 14590
rect 207150 14520 207350 14590
rect 207650 14520 207850 14590
rect 204150 14410 204350 14480
rect 204650 14410 204850 14480
rect 205150 14410 205350 14480
rect 205650 14410 205850 14480
rect 206150 14410 206350 14480
rect 206650 14410 206850 14480
rect 207150 14410 207350 14480
rect 207650 14410 207850 14480
rect 204020 14150 204090 14350
rect 204410 14150 204480 14350
rect 204520 14150 204590 14350
rect 204910 14150 204980 14350
rect 205020 14150 205090 14350
rect 205410 14150 205480 14350
rect 205520 14150 205590 14350
rect 205910 14150 205980 14350
rect 206020 14150 206090 14350
rect 206410 14150 206480 14350
rect 206520 14150 206590 14350
rect 206910 14150 206980 14350
rect 207020 14150 207090 14350
rect 207410 14150 207480 14350
rect 207520 14150 207590 14350
rect 207910 14150 207980 14350
rect 204150 14020 204350 14090
rect 204650 14020 204850 14090
rect 205150 14020 205350 14090
rect 205650 14020 205850 14090
rect 206150 14020 206350 14090
rect 206650 14020 206850 14090
rect 207150 14020 207350 14090
rect 207650 14020 207850 14090
rect 204150 13910 204350 13980
rect 204650 13910 204850 13980
rect 205150 13910 205350 13980
rect 205650 13910 205850 13980
rect 206150 13910 206350 13980
rect 206650 13910 206850 13980
rect 207150 13910 207350 13980
rect 207650 13910 207850 13980
rect 204020 13650 204090 13850
rect 204410 13650 204480 13850
rect 204520 13650 204590 13850
rect 204910 13650 204980 13850
rect 205020 13650 205090 13850
rect 205410 13650 205480 13850
rect 205520 13650 205590 13850
rect 205910 13650 205980 13850
rect 206020 13650 206090 13850
rect 206410 13650 206480 13850
rect 206520 13650 206590 13850
rect 206910 13650 206980 13850
rect 207020 13650 207090 13850
rect 207410 13650 207480 13850
rect 207520 13650 207590 13850
rect 207910 13650 207980 13850
rect 204150 13520 204350 13590
rect 204650 13520 204850 13590
rect 205150 13520 205350 13590
rect 205650 13520 205850 13590
rect 206150 13520 206350 13590
rect 206650 13520 206850 13590
rect 207150 13520 207350 13590
rect 207650 13520 207850 13590
rect 204150 13410 204350 13480
rect 204650 13410 204850 13480
rect 205150 13410 205350 13480
rect 205650 13410 205850 13480
rect 206150 13410 206350 13480
rect 206650 13410 206850 13480
rect 207150 13410 207350 13480
rect 207650 13410 207850 13480
rect 204020 13150 204090 13350
rect 204410 13150 204480 13350
rect 204520 13150 204590 13350
rect 204910 13150 204980 13350
rect 205020 13150 205090 13350
rect 205410 13150 205480 13350
rect 205520 13150 205590 13350
rect 205910 13150 205980 13350
rect 206020 13150 206090 13350
rect 206410 13150 206480 13350
rect 206520 13150 206590 13350
rect 206910 13150 206980 13350
rect 207020 13150 207090 13350
rect 207410 13150 207480 13350
rect 207520 13150 207590 13350
rect 207910 13150 207980 13350
rect 204150 13020 204350 13090
rect 204650 13020 204850 13090
rect 205150 13020 205350 13090
rect 205650 13020 205850 13090
rect 206150 13020 206350 13090
rect 206650 13020 206850 13090
rect 207150 13020 207350 13090
rect 207650 13020 207850 13090
rect 204150 12910 204350 12980
rect 204650 12910 204850 12980
rect 205150 12910 205350 12980
rect 205650 12910 205850 12980
rect 206150 12910 206350 12980
rect 206650 12910 206850 12980
rect 207150 12910 207350 12980
rect 207650 12910 207850 12980
rect 204020 12650 204090 12850
rect 204410 12650 204480 12850
rect 204520 12650 204590 12850
rect 204910 12650 204980 12850
rect 205020 12650 205090 12850
rect 205410 12650 205480 12850
rect 205520 12650 205590 12850
rect 205910 12650 205980 12850
rect 206020 12650 206090 12850
rect 206410 12650 206480 12850
rect 206520 12650 206590 12850
rect 206910 12650 206980 12850
rect 207020 12650 207090 12850
rect 207410 12650 207480 12850
rect 207520 12650 207590 12850
rect 207910 12650 207980 12850
rect 204150 12520 204350 12590
rect 204650 12520 204850 12590
rect 205150 12520 205350 12590
rect 205650 12520 205850 12590
rect 206150 12520 206350 12590
rect 206650 12520 206850 12590
rect 207150 12520 207350 12590
rect 207650 12520 207850 12590
rect 204150 12410 204350 12480
rect 204650 12410 204850 12480
rect 205150 12410 205350 12480
rect 205650 12410 205850 12480
rect 206150 12410 206350 12480
rect 206650 12410 206850 12480
rect 207150 12410 207350 12480
rect 207650 12410 207850 12480
rect 204020 12150 204090 12350
rect 204410 12150 204480 12350
rect 204520 12150 204590 12350
rect 204910 12150 204980 12350
rect 205020 12150 205090 12350
rect 205410 12150 205480 12350
rect 205520 12150 205590 12350
rect 205910 12150 205980 12350
rect 206020 12150 206090 12350
rect 206410 12150 206480 12350
rect 206520 12150 206590 12350
rect 206910 12150 206980 12350
rect 207020 12150 207090 12350
rect 207410 12150 207480 12350
rect 207520 12150 207590 12350
rect 207910 12150 207980 12350
rect 204150 12020 204350 12090
rect 204650 12020 204850 12090
rect 205150 12020 205350 12090
rect 205650 12020 205850 12090
rect 206150 12020 206350 12090
rect 206650 12020 206850 12090
rect 207150 12020 207350 12090
rect 207650 12020 207850 12090
rect 204150 11910 204350 11980
rect 204650 11910 204850 11980
rect 205150 11910 205350 11980
rect 205650 11910 205850 11980
rect 206150 11910 206350 11980
rect 206650 11910 206850 11980
rect 207150 11910 207350 11980
rect 207650 11910 207850 11980
rect 204020 11650 204090 11850
rect 204410 11650 204480 11850
rect 204520 11650 204590 11850
rect 204910 11650 204980 11850
rect 205020 11650 205090 11850
rect 205410 11650 205480 11850
rect 205520 11650 205590 11850
rect 205910 11650 205980 11850
rect 206020 11650 206090 11850
rect 206410 11650 206480 11850
rect 206520 11650 206590 11850
rect 206910 11650 206980 11850
rect 207020 11650 207090 11850
rect 207410 11650 207480 11850
rect 207520 11650 207590 11850
rect 207910 11650 207980 11850
rect 204150 11520 204350 11590
rect 204650 11520 204850 11590
rect 205150 11520 205350 11590
rect 205650 11520 205850 11590
rect 206150 11520 206350 11590
rect 206650 11520 206850 11590
rect 207150 11520 207350 11590
rect 207650 11520 207850 11590
rect 204150 11410 204350 11480
rect 204650 11410 204850 11480
rect 205150 11410 205350 11480
rect 205650 11410 205850 11480
rect 206150 11410 206350 11480
rect 206650 11410 206850 11480
rect 207150 11410 207350 11480
rect 207650 11410 207850 11480
rect 204020 11150 204090 11350
rect 204410 11150 204480 11350
rect 204520 11150 204590 11350
rect 204910 11150 204980 11350
rect 205020 11150 205090 11350
rect 205410 11150 205480 11350
rect 205520 11150 205590 11350
rect 205910 11150 205980 11350
rect 206020 11150 206090 11350
rect 206410 11150 206480 11350
rect 206520 11150 206590 11350
rect 206910 11150 206980 11350
rect 207020 11150 207090 11350
rect 207410 11150 207480 11350
rect 207520 11150 207590 11350
rect 207910 11150 207980 11350
rect 204150 11020 204350 11090
rect 204650 11020 204850 11090
rect 205150 11020 205350 11090
rect 205650 11020 205850 11090
rect 206150 11020 206350 11090
rect 206650 11020 206850 11090
rect 207150 11020 207350 11090
rect 207650 11020 207850 11090
rect 204150 10910 204350 10980
rect 204650 10910 204850 10980
rect 205150 10910 205350 10980
rect 205650 10910 205850 10980
rect 206150 10910 206350 10980
rect 206650 10910 206850 10980
rect 207150 10910 207350 10980
rect 207650 10910 207850 10980
rect 204020 10650 204090 10850
rect 204410 10650 204480 10850
rect 204520 10650 204590 10850
rect 204910 10650 204980 10850
rect 205020 10650 205090 10850
rect 205410 10650 205480 10850
rect 205520 10650 205590 10850
rect 205910 10650 205980 10850
rect 206020 10650 206090 10850
rect 206410 10650 206480 10850
rect 206520 10650 206590 10850
rect 206910 10650 206980 10850
rect 207020 10650 207090 10850
rect 207410 10650 207480 10850
rect 207520 10650 207590 10850
rect 207910 10650 207980 10850
rect 204150 10520 204350 10590
rect 204650 10520 204850 10590
rect 205150 10520 205350 10590
rect 205650 10520 205850 10590
rect 206150 10520 206350 10590
rect 206650 10520 206850 10590
rect 207150 10520 207350 10590
rect 207650 10520 207850 10590
rect 204150 10410 204350 10480
rect 204650 10410 204850 10480
rect 205150 10410 205350 10480
rect 205650 10410 205850 10480
rect 206150 10410 206350 10480
rect 206650 10410 206850 10480
rect 207150 10410 207350 10480
rect 207650 10410 207850 10480
rect 204020 10150 204090 10350
rect 204410 10150 204480 10350
rect 204520 10150 204590 10350
rect 204910 10150 204980 10350
rect 205020 10150 205090 10350
rect 205410 10150 205480 10350
rect 205520 10150 205590 10350
rect 205910 10150 205980 10350
rect 206020 10150 206090 10350
rect 206410 10150 206480 10350
rect 206520 10150 206590 10350
rect 206910 10150 206980 10350
rect 207020 10150 207090 10350
rect 207410 10150 207480 10350
rect 207520 10150 207590 10350
rect 207910 10150 207980 10350
rect 204150 10020 204350 10090
rect 204650 10020 204850 10090
rect 205150 10020 205350 10090
rect 205650 10020 205850 10090
rect 206150 10020 206350 10090
rect 206650 10020 206850 10090
rect 207150 10020 207350 10090
rect 207650 10020 207850 10090
rect 204150 9910 204350 9980
rect 204650 9910 204850 9980
rect 205150 9910 205350 9980
rect 205650 9910 205850 9980
rect 206150 9910 206350 9980
rect 206650 9910 206850 9980
rect 207150 9910 207350 9980
rect 207650 9910 207850 9980
rect 204020 9650 204090 9850
rect 204410 9650 204480 9850
rect 204520 9650 204590 9850
rect 204910 9650 204980 9850
rect 205020 9650 205090 9850
rect 205410 9650 205480 9850
rect 205520 9650 205590 9850
rect 205910 9650 205980 9850
rect 206020 9650 206090 9850
rect 206410 9650 206480 9850
rect 206520 9650 206590 9850
rect 206910 9650 206980 9850
rect 207020 9650 207090 9850
rect 207410 9650 207480 9850
rect 207520 9650 207590 9850
rect 207910 9650 207980 9850
rect 204150 9520 204350 9590
rect 204650 9520 204850 9590
rect 205150 9520 205350 9590
rect 205650 9520 205850 9590
rect 206150 9520 206350 9590
rect 206650 9520 206850 9590
rect 207150 9520 207350 9590
rect 207650 9520 207850 9590
rect 204150 9410 204350 9480
rect 204650 9410 204850 9480
rect 205150 9410 205350 9480
rect 205650 9410 205850 9480
rect 206150 9410 206350 9480
rect 206650 9410 206850 9480
rect 207150 9410 207350 9480
rect 207650 9410 207850 9480
rect 204020 9150 204090 9350
rect 204410 9150 204480 9350
rect 204520 9150 204590 9350
rect 204910 9150 204980 9350
rect 205020 9150 205090 9350
rect 205410 9150 205480 9350
rect 205520 9150 205590 9350
rect 205910 9150 205980 9350
rect 206020 9150 206090 9350
rect 206410 9150 206480 9350
rect 206520 9150 206590 9350
rect 206910 9150 206980 9350
rect 207020 9150 207090 9350
rect 207410 9150 207480 9350
rect 207520 9150 207590 9350
rect 207910 9150 207980 9350
rect 204150 9020 204350 9090
rect 204650 9020 204850 9090
rect 205150 9020 205350 9090
rect 205650 9020 205850 9090
rect 206150 9020 206350 9090
rect 206650 9020 206850 9090
rect 207150 9020 207350 9090
rect 207650 9020 207850 9090
rect 204150 8910 204350 8980
rect 204650 8910 204850 8980
rect 205150 8910 205350 8980
rect 205650 8910 205850 8980
rect 206150 8910 206350 8980
rect 206650 8910 206850 8980
rect 207150 8910 207350 8980
rect 207650 8910 207850 8980
rect 204020 8650 204090 8850
rect 204410 8650 204480 8850
rect 204520 8650 204590 8850
rect 204910 8650 204980 8850
rect 205020 8650 205090 8850
rect 205410 8650 205480 8850
rect 205520 8650 205590 8850
rect 205910 8650 205980 8850
rect 206020 8650 206090 8850
rect 206410 8650 206480 8850
rect 206520 8650 206590 8850
rect 206910 8650 206980 8850
rect 207020 8650 207090 8850
rect 207410 8650 207480 8850
rect 207520 8650 207590 8850
rect 207910 8650 207980 8850
rect 204150 8520 204350 8590
rect 204650 8520 204850 8590
rect 205150 8520 205350 8590
rect 205650 8520 205850 8590
rect 206150 8520 206350 8590
rect 206650 8520 206850 8590
rect 207150 8520 207350 8590
rect 207650 8520 207850 8590
rect 204150 8410 204350 8480
rect 204650 8410 204850 8480
rect 205150 8410 205350 8480
rect 205650 8410 205850 8480
rect 206150 8410 206350 8480
rect 206650 8410 206850 8480
rect 207150 8410 207350 8480
rect 207650 8410 207850 8480
rect 204020 8150 204090 8350
rect 204410 8150 204480 8350
rect 204520 8150 204590 8350
rect 204910 8150 204980 8350
rect 205020 8150 205090 8350
rect 205410 8150 205480 8350
rect 205520 8150 205590 8350
rect 205910 8150 205980 8350
rect 206020 8150 206090 8350
rect 206410 8150 206480 8350
rect 206520 8150 206590 8350
rect 206910 8150 206980 8350
rect 207020 8150 207090 8350
rect 207410 8150 207480 8350
rect 207520 8150 207590 8350
rect 207910 8150 207980 8350
rect 204150 8020 204350 8090
rect 204650 8020 204850 8090
rect 205150 8020 205350 8090
rect 205650 8020 205850 8090
rect 206150 8020 206350 8090
rect 206650 8020 206850 8090
rect 207150 8020 207350 8090
rect 207650 8020 207850 8090
rect 204150 7910 204350 7980
rect 204650 7910 204850 7980
rect 205150 7910 205350 7980
rect 205650 7910 205850 7980
rect 206150 7910 206350 7980
rect 206650 7910 206850 7980
rect 207150 7910 207350 7980
rect 207650 7910 207850 7980
rect 204020 7650 204090 7850
rect 204410 7650 204480 7850
rect 204520 7650 204590 7850
rect 204910 7650 204980 7850
rect 205020 7650 205090 7850
rect 205410 7650 205480 7850
rect 205520 7650 205590 7850
rect 205910 7650 205980 7850
rect 206020 7650 206090 7850
rect 206410 7650 206480 7850
rect 206520 7650 206590 7850
rect 206910 7650 206980 7850
rect 207020 7650 207090 7850
rect 207410 7650 207480 7850
rect 207520 7650 207590 7850
rect 207910 7650 207980 7850
rect 204150 7520 204350 7590
rect 204650 7520 204850 7590
rect 205150 7520 205350 7590
rect 205650 7520 205850 7590
rect 206150 7520 206350 7590
rect 206650 7520 206850 7590
rect 207150 7520 207350 7590
rect 207650 7520 207850 7590
rect 204150 7410 204350 7480
rect 204650 7410 204850 7480
rect 205150 7410 205350 7480
rect 205650 7410 205850 7480
rect 206150 7410 206350 7480
rect 206650 7410 206850 7480
rect 207150 7410 207350 7480
rect 207650 7410 207850 7480
rect 204020 7150 204090 7350
rect 204410 7150 204480 7350
rect 204520 7150 204590 7350
rect 204910 7150 204980 7350
rect 205020 7150 205090 7350
rect 205410 7150 205480 7350
rect 205520 7150 205590 7350
rect 205910 7150 205980 7350
rect 206020 7150 206090 7350
rect 206410 7150 206480 7350
rect 206520 7150 206590 7350
rect 206910 7150 206980 7350
rect 207020 7150 207090 7350
rect 207410 7150 207480 7350
rect 207520 7150 207590 7350
rect 207910 7150 207980 7350
rect 204150 7020 204350 7090
rect 204650 7020 204850 7090
rect 205150 7020 205350 7090
rect 205650 7020 205850 7090
rect 206150 7020 206350 7090
rect 206650 7020 206850 7090
rect 207150 7020 207350 7090
rect 207650 7020 207850 7090
rect 204150 6910 204350 6980
rect 204650 6910 204850 6980
rect 205150 6910 205350 6980
rect 205650 6910 205850 6980
rect 206150 6910 206350 6980
rect 206650 6910 206850 6980
rect 207150 6910 207350 6980
rect 207650 6910 207850 6980
rect 204020 6650 204090 6850
rect 204410 6650 204480 6850
rect 204520 6650 204590 6850
rect 204910 6650 204980 6850
rect 205020 6650 205090 6850
rect 205410 6650 205480 6850
rect 205520 6650 205590 6850
rect 205910 6650 205980 6850
rect 206020 6650 206090 6850
rect 206410 6650 206480 6850
rect 206520 6650 206590 6850
rect 206910 6650 206980 6850
rect 207020 6650 207090 6850
rect 207410 6650 207480 6850
rect 207520 6650 207590 6850
rect 207910 6650 207980 6850
rect 204150 6520 204350 6590
rect 204650 6520 204850 6590
rect 205150 6520 205350 6590
rect 205650 6520 205850 6590
rect 206150 6520 206350 6590
rect 206650 6520 206850 6590
rect 207150 6520 207350 6590
rect 207650 6520 207850 6590
rect 204150 6410 204350 6480
rect 204650 6410 204850 6480
rect 205150 6410 205350 6480
rect 205650 6410 205850 6480
rect 206150 6410 206350 6480
rect 206650 6410 206850 6480
rect 207150 6410 207350 6480
rect 207650 6410 207850 6480
rect 204020 6150 204090 6350
rect 204410 6150 204480 6350
rect 204520 6150 204590 6350
rect 204910 6150 204980 6350
rect 205020 6150 205090 6350
rect 205410 6150 205480 6350
rect 205520 6150 205590 6350
rect 205910 6150 205980 6350
rect 206020 6150 206090 6350
rect 206410 6150 206480 6350
rect 206520 6150 206590 6350
rect 206910 6150 206980 6350
rect 207020 6150 207090 6350
rect 207410 6150 207480 6350
rect 207520 6150 207590 6350
rect 207910 6150 207980 6350
rect 204150 6020 204350 6090
rect 204650 6020 204850 6090
rect 205150 6020 205350 6090
rect 205650 6020 205850 6090
rect 206150 6020 206350 6090
rect 206650 6020 206850 6090
rect 207150 6020 207350 6090
rect 207650 6020 207850 6090
rect 198150 5910 198350 5980
rect 198650 5910 198850 5980
rect 199150 5910 199350 5980
rect 199650 5910 199850 5980
rect 200150 5910 200350 5980
rect 200650 5910 200850 5980
rect 201150 5910 201350 5980
rect 201650 5910 201850 5980
rect 202150 5910 202350 5980
rect 202650 5910 202850 5980
rect 203150 5910 203350 5980
rect 203650 5910 203850 5980
rect 204150 5910 204350 5980
rect 204650 5910 204850 5980
rect 205150 5910 205350 5980
rect 205650 5910 205850 5980
rect 206150 5910 206350 5980
rect 206650 5910 206850 5980
rect 207150 5910 207350 5980
rect 207650 5910 207850 5980
rect 198020 5650 198090 5850
rect 198410 5650 198480 5850
rect 198520 5650 198590 5850
rect 198910 5650 198980 5850
rect 199020 5650 199090 5850
rect 199410 5650 199480 5850
rect 199520 5650 199590 5850
rect 199910 5650 199980 5850
rect 200020 5650 200090 5850
rect 200410 5650 200480 5850
rect 200520 5650 200590 5850
rect 200910 5650 200980 5850
rect 201020 5650 201090 5850
rect 201410 5650 201480 5850
rect 201520 5650 201590 5850
rect 201910 5650 201980 5850
rect 202020 5650 202090 5850
rect 202410 5650 202480 5850
rect 202520 5650 202590 5850
rect 202910 5650 202980 5850
rect 203020 5650 203090 5850
rect 203410 5650 203480 5850
rect 203520 5650 203590 5850
rect 203910 5650 203980 5850
rect 204020 5650 204090 5850
rect 204410 5650 204480 5850
rect 204520 5650 204590 5850
rect 204910 5650 204980 5850
rect 205020 5650 205090 5850
rect 205410 5650 205480 5850
rect 205520 5650 205590 5850
rect 205910 5650 205980 5850
rect 206020 5650 206090 5850
rect 206410 5650 206480 5850
rect 206520 5650 206590 5850
rect 206910 5650 206980 5850
rect 207020 5650 207090 5850
rect 207410 5650 207480 5850
rect 207520 5650 207590 5850
rect 207910 5650 207980 5850
rect 198150 5520 198350 5590
rect 198650 5520 198850 5590
rect 199150 5520 199350 5590
rect 199650 5520 199850 5590
rect 200150 5520 200350 5590
rect 200650 5520 200850 5590
rect 201150 5520 201350 5590
rect 201650 5520 201850 5590
rect 202150 5520 202350 5590
rect 202650 5520 202850 5590
rect 203150 5520 203350 5590
rect 203650 5520 203850 5590
rect 204150 5520 204350 5590
rect 204650 5520 204850 5590
rect 205150 5520 205350 5590
rect 205650 5520 205850 5590
rect 206150 5520 206350 5590
rect 206650 5520 206850 5590
rect 207150 5520 207350 5590
rect 207650 5520 207850 5590
rect 198150 5410 198350 5480
rect 198650 5410 198850 5480
rect 199150 5410 199350 5480
rect 199650 5410 199850 5480
rect 200150 5410 200350 5480
rect 200650 5410 200850 5480
rect 201150 5410 201350 5480
rect 201650 5410 201850 5480
rect 202150 5410 202350 5480
rect 202650 5410 202850 5480
rect 203150 5410 203350 5480
rect 203650 5410 203850 5480
rect 204150 5410 204350 5480
rect 204650 5410 204850 5480
rect 205150 5410 205350 5480
rect 205650 5410 205850 5480
rect 206150 5410 206350 5480
rect 206650 5410 206850 5480
rect 207150 5410 207350 5480
rect 207650 5410 207850 5480
rect 198020 5150 198090 5350
rect 198410 5150 198480 5350
rect 198520 5150 198590 5350
rect 198910 5150 198980 5350
rect 199020 5150 199090 5350
rect 199410 5150 199480 5350
rect 199520 5150 199590 5350
rect 199910 5150 199980 5350
rect 200020 5150 200090 5350
rect 200410 5150 200480 5350
rect 200520 5150 200590 5350
rect 200910 5150 200980 5350
rect 201020 5150 201090 5350
rect 201410 5150 201480 5350
rect 201520 5150 201590 5350
rect 201910 5150 201980 5350
rect 202020 5150 202090 5350
rect 202410 5150 202480 5350
rect 202520 5150 202590 5350
rect 202910 5150 202980 5350
rect 203020 5150 203090 5350
rect 203410 5150 203480 5350
rect 203520 5150 203590 5350
rect 203910 5150 203980 5350
rect 204020 5150 204090 5350
rect 204410 5150 204480 5350
rect 204520 5150 204590 5350
rect 204910 5150 204980 5350
rect 205020 5150 205090 5350
rect 205410 5150 205480 5350
rect 205520 5150 205590 5350
rect 205910 5150 205980 5350
rect 206020 5150 206090 5350
rect 206410 5150 206480 5350
rect 206520 5150 206590 5350
rect 206910 5150 206980 5350
rect 207020 5150 207090 5350
rect 207410 5150 207480 5350
rect 207520 5150 207590 5350
rect 207910 5150 207980 5350
rect 198150 5020 198350 5090
rect 198650 5020 198850 5090
rect 199150 5020 199350 5090
rect 199650 5020 199850 5090
rect 200150 5020 200350 5090
rect 200650 5020 200850 5090
rect 201150 5020 201350 5090
rect 201650 5020 201850 5090
rect 202150 5020 202350 5090
rect 202650 5020 202850 5090
rect 203150 5020 203350 5090
rect 203650 5020 203850 5090
rect 204150 5020 204350 5090
rect 204650 5020 204850 5090
rect 205150 5020 205350 5090
rect 205650 5020 205850 5090
rect 206150 5020 206350 5090
rect 206650 5020 206850 5090
rect 207150 5020 207350 5090
rect 207650 5020 207850 5090
rect 198150 4910 198350 4980
rect 198650 4910 198850 4980
rect 199150 4910 199350 4980
rect 199650 4910 199850 4980
rect 200150 4910 200350 4980
rect 200650 4910 200850 4980
rect 201150 4910 201350 4980
rect 201650 4910 201850 4980
rect 202150 4910 202350 4980
rect 202650 4910 202850 4980
rect 203150 4910 203350 4980
rect 203650 4910 203850 4980
rect 204150 4910 204350 4980
rect 204650 4910 204850 4980
rect 205150 4910 205350 4980
rect 205650 4910 205850 4980
rect 206150 4910 206350 4980
rect 206650 4910 206850 4980
rect 207150 4910 207350 4980
rect 207650 4910 207850 4980
rect 198020 4650 198090 4850
rect 198410 4650 198480 4850
rect 198520 4650 198590 4850
rect 198910 4650 198980 4850
rect 199020 4650 199090 4850
rect 199410 4650 199480 4850
rect 199520 4650 199590 4850
rect 199910 4650 199980 4850
rect 200020 4650 200090 4850
rect 200410 4650 200480 4850
rect 200520 4650 200590 4850
rect 200910 4650 200980 4850
rect 201020 4650 201090 4850
rect 201410 4650 201480 4850
rect 201520 4650 201590 4850
rect 201910 4650 201980 4850
rect 202020 4650 202090 4850
rect 202410 4650 202480 4850
rect 202520 4650 202590 4850
rect 202910 4650 202980 4850
rect 203020 4650 203090 4850
rect 203410 4650 203480 4850
rect 203520 4650 203590 4850
rect 203910 4650 203980 4850
rect 204020 4650 204090 4850
rect 204410 4650 204480 4850
rect 204520 4650 204590 4850
rect 204910 4650 204980 4850
rect 205020 4650 205090 4850
rect 205410 4650 205480 4850
rect 205520 4650 205590 4850
rect 205910 4650 205980 4850
rect 206020 4650 206090 4850
rect 206410 4650 206480 4850
rect 206520 4650 206590 4850
rect 206910 4650 206980 4850
rect 207020 4650 207090 4850
rect 207410 4650 207480 4850
rect 207520 4650 207590 4850
rect 207910 4650 207980 4850
rect 198150 4520 198350 4590
rect 198650 4520 198850 4590
rect 199150 4520 199350 4590
rect 199650 4520 199850 4590
rect 200150 4520 200350 4590
rect 200650 4520 200850 4590
rect 201150 4520 201350 4590
rect 201650 4520 201850 4590
rect 202150 4520 202350 4590
rect 202650 4520 202850 4590
rect 203150 4520 203350 4590
rect 203650 4520 203850 4590
rect 204150 4520 204350 4590
rect 204650 4520 204850 4590
rect 205150 4520 205350 4590
rect 205650 4520 205850 4590
rect 206150 4520 206350 4590
rect 206650 4520 206850 4590
rect 207150 4520 207350 4590
rect 207650 4520 207850 4590
rect 198150 4410 198350 4480
rect 198650 4410 198850 4480
rect 199150 4410 199350 4480
rect 199650 4410 199850 4480
rect 200150 4410 200350 4480
rect 200650 4410 200850 4480
rect 201150 4410 201350 4480
rect 201650 4410 201850 4480
rect 202150 4410 202350 4480
rect 202650 4410 202850 4480
rect 203150 4410 203350 4480
rect 203650 4410 203850 4480
rect 204150 4410 204350 4480
rect 204650 4410 204850 4480
rect 205150 4410 205350 4480
rect 205650 4410 205850 4480
rect 206150 4410 206350 4480
rect 206650 4410 206850 4480
rect 207150 4410 207350 4480
rect 207650 4410 207850 4480
rect 198020 4150 198090 4350
rect 198410 4150 198480 4350
rect 198520 4150 198590 4350
rect 198910 4150 198980 4350
rect 199020 4150 199090 4350
rect 199410 4150 199480 4350
rect 199520 4150 199590 4350
rect 199910 4150 199980 4350
rect 200020 4150 200090 4350
rect 200410 4150 200480 4350
rect 200520 4150 200590 4350
rect 200910 4150 200980 4350
rect 201020 4150 201090 4350
rect 201410 4150 201480 4350
rect 201520 4150 201590 4350
rect 201910 4150 201980 4350
rect 202020 4150 202090 4350
rect 202410 4150 202480 4350
rect 202520 4150 202590 4350
rect 202910 4150 202980 4350
rect 203020 4150 203090 4350
rect 203410 4150 203480 4350
rect 203520 4150 203590 4350
rect 203910 4150 203980 4350
rect 204020 4150 204090 4350
rect 204410 4150 204480 4350
rect 204520 4150 204590 4350
rect 204910 4150 204980 4350
rect 205020 4150 205090 4350
rect 205410 4150 205480 4350
rect 205520 4150 205590 4350
rect 205910 4150 205980 4350
rect 206020 4150 206090 4350
rect 206410 4150 206480 4350
rect 206520 4150 206590 4350
rect 206910 4150 206980 4350
rect 207020 4150 207090 4350
rect 207410 4150 207480 4350
rect 207520 4150 207590 4350
rect 207910 4150 207980 4350
rect 198150 4020 198350 4090
rect 198650 4020 198850 4090
rect 199150 4020 199350 4090
rect 199650 4020 199850 4090
rect 200150 4020 200350 4090
rect 200650 4020 200850 4090
rect 201150 4020 201350 4090
rect 201650 4020 201850 4090
rect 202150 4020 202350 4090
rect 202650 4020 202850 4090
rect 203150 4020 203350 4090
rect 203650 4020 203850 4090
rect 204150 4020 204350 4090
rect 204650 4020 204850 4090
rect 205150 4020 205350 4090
rect 205650 4020 205850 4090
rect 206150 4020 206350 4090
rect 206650 4020 206850 4090
rect 207150 4020 207350 4090
rect 207650 4020 207850 4090
rect 198150 3910 198350 3980
rect 198650 3910 198850 3980
rect 199150 3910 199350 3980
rect 199650 3910 199850 3980
rect 200150 3910 200350 3980
rect 200650 3910 200850 3980
rect 201150 3910 201350 3980
rect 201650 3910 201850 3980
rect 202150 3910 202350 3980
rect 202650 3910 202850 3980
rect 203150 3910 203350 3980
rect 203650 3910 203850 3980
rect 204150 3910 204350 3980
rect 204650 3910 204850 3980
rect 205150 3910 205350 3980
rect 205650 3910 205850 3980
rect 206150 3910 206350 3980
rect 206650 3910 206850 3980
rect 207150 3910 207350 3980
rect 207650 3910 207850 3980
rect 198020 3650 198090 3850
rect 198410 3650 198480 3850
rect 198520 3650 198590 3850
rect 198910 3650 198980 3850
rect 199020 3650 199090 3850
rect 199410 3650 199480 3850
rect 199520 3650 199590 3850
rect 199910 3650 199980 3850
rect 200020 3650 200090 3850
rect 200410 3650 200480 3850
rect 200520 3650 200590 3850
rect 200910 3650 200980 3850
rect 201020 3650 201090 3850
rect 201410 3650 201480 3850
rect 201520 3650 201590 3850
rect 201910 3650 201980 3850
rect 202020 3650 202090 3850
rect 202410 3650 202480 3850
rect 202520 3650 202590 3850
rect 202910 3650 202980 3850
rect 203020 3650 203090 3850
rect 203410 3650 203480 3850
rect 203520 3650 203590 3850
rect 203910 3650 203980 3850
rect 204020 3650 204090 3850
rect 204410 3650 204480 3850
rect 204520 3650 204590 3850
rect 204910 3650 204980 3850
rect 205020 3650 205090 3850
rect 205410 3650 205480 3850
rect 205520 3650 205590 3850
rect 205910 3650 205980 3850
rect 206020 3650 206090 3850
rect 206410 3650 206480 3850
rect 206520 3650 206590 3850
rect 206910 3650 206980 3850
rect 207020 3650 207090 3850
rect 207410 3650 207480 3850
rect 207520 3650 207590 3850
rect 207910 3650 207980 3850
rect 198150 3520 198350 3590
rect 198650 3520 198850 3590
rect 199150 3520 199350 3590
rect 199650 3520 199850 3590
rect 200150 3520 200350 3590
rect 200650 3520 200850 3590
rect 201150 3520 201350 3590
rect 201650 3520 201850 3590
rect 202150 3520 202350 3590
rect 202650 3520 202850 3590
rect 203150 3520 203350 3590
rect 203650 3520 203850 3590
rect 204150 3520 204350 3590
rect 204650 3520 204850 3590
rect 205150 3520 205350 3590
rect 205650 3520 205850 3590
rect 206150 3520 206350 3590
rect 206650 3520 206850 3590
rect 207150 3520 207350 3590
rect 207650 3520 207850 3590
rect 198150 3410 198350 3480
rect 198650 3410 198850 3480
rect 199150 3410 199350 3480
rect 199650 3410 199850 3480
rect 200150 3410 200350 3480
rect 200650 3410 200850 3480
rect 201150 3410 201350 3480
rect 201650 3410 201850 3480
rect 202150 3410 202350 3480
rect 202650 3410 202850 3480
rect 203150 3410 203350 3480
rect 203650 3410 203850 3480
rect 204150 3410 204350 3480
rect 204650 3410 204850 3480
rect 205150 3410 205350 3480
rect 205650 3410 205850 3480
rect 206150 3410 206350 3480
rect 206650 3410 206850 3480
rect 207150 3410 207350 3480
rect 207650 3410 207850 3480
rect 198020 3150 198090 3350
rect 198410 3150 198480 3350
rect 198520 3150 198590 3350
rect 198910 3150 198980 3350
rect 199020 3150 199090 3350
rect 199410 3150 199480 3350
rect 199520 3150 199590 3350
rect 199910 3150 199980 3350
rect 200020 3150 200090 3350
rect 200410 3150 200480 3350
rect 200520 3150 200590 3350
rect 200910 3150 200980 3350
rect 201020 3150 201090 3350
rect 201410 3150 201480 3350
rect 201520 3150 201590 3350
rect 201910 3150 201980 3350
rect 202020 3150 202090 3350
rect 202410 3150 202480 3350
rect 202520 3150 202590 3350
rect 202910 3150 202980 3350
rect 203020 3150 203090 3350
rect 203410 3150 203480 3350
rect 203520 3150 203590 3350
rect 203910 3150 203980 3350
rect 204020 3150 204090 3350
rect 204410 3150 204480 3350
rect 204520 3150 204590 3350
rect 204910 3150 204980 3350
rect 205020 3150 205090 3350
rect 205410 3150 205480 3350
rect 205520 3150 205590 3350
rect 205910 3150 205980 3350
rect 206020 3150 206090 3350
rect 206410 3150 206480 3350
rect 206520 3150 206590 3350
rect 206910 3150 206980 3350
rect 207020 3150 207090 3350
rect 207410 3150 207480 3350
rect 207520 3150 207590 3350
rect 207910 3150 207980 3350
rect 198150 3020 198350 3090
rect 198650 3020 198850 3090
rect 199150 3020 199350 3090
rect 199650 3020 199850 3090
rect 200150 3020 200350 3090
rect 200650 3020 200850 3090
rect 201150 3020 201350 3090
rect 201650 3020 201850 3090
rect 202150 3020 202350 3090
rect 202650 3020 202850 3090
rect 203150 3020 203350 3090
rect 203650 3020 203850 3090
rect 204150 3020 204350 3090
rect 204650 3020 204850 3090
rect 205150 3020 205350 3090
rect 205650 3020 205850 3090
rect 206150 3020 206350 3090
rect 206650 3020 206850 3090
rect 207150 3020 207350 3090
rect 207650 3020 207850 3090
rect 198150 2910 198350 2980
rect 198650 2910 198850 2980
rect 199150 2910 199350 2980
rect 199650 2910 199850 2980
rect 200150 2910 200350 2980
rect 200650 2910 200850 2980
rect 201150 2910 201350 2980
rect 201650 2910 201850 2980
rect 202150 2910 202350 2980
rect 202650 2910 202850 2980
rect 203150 2910 203350 2980
rect 203650 2910 203850 2980
rect 204150 2910 204350 2980
rect 204650 2910 204850 2980
rect 205150 2910 205350 2980
rect 205650 2910 205850 2980
rect 206150 2910 206350 2980
rect 206650 2910 206850 2980
rect 207150 2910 207350 2980
rect 207650 2910 207850 2980
rect 198020 2650 198090 2850
rect 198410 2650 198480 2850
rect 198520 2650 198590 2850
rect 198910 2650 198980 2850
rect 199020 2650 199090 2850
rect 199410 2650 199480 2850
rect 199520 2650 199590 2850
rect 199910 2650 199980 2850
rect 200020 2650 200090 2850
rect 200410 2650 200480 2850
rect 200520 2650 200590 2850
rect 200910 2650 200980 2850
rect 201020 2650 201090 2850
rect 201410 2650 201480 2850
rect 201520 2650 201590 2850
rect 201910 2650 201980 2850
rect 202020 2650 202090 2850
rect 202410 2650 202480 2850
rect 202520 2650 202590 2850
rect 202910 2650 202980 2850
rect 203020 2650 203090 2850
rect 203410 2650 203480 2850
rect 203520 2650 203590 2850
rect 203910 2650 203980 2850
rect 204020 2650 204090 2850
rect 204410 2650 204480 2850
rect 204520 2650 204590 2850
rect 204910 2650 204980 2850
rect 205020 2650 205090 2850
rect 205410 2650 205480 2850
rect 205520 2650 205590 2850
rect 205910 2650 205980 2850
rect 206020 2650 206090 2850
rect 206410 2650 206480 2850
rect 206520 2650 206590 2850
rect 206910 2650 206980 2850
rect 207020 2650 207090 2850
rect 207410 2650 207480 2850
rect 207520 2650 207590 2850
rect 207910 2650 207980 2850
rect 198150 2520 198350 2590
rect 198650 2520 198850 2590
rect 199150 2520 199350 2590
rect 199650 2520 199850 2590
rect 200150 2520 200350 2590
rect 200650 2520 200850 2590
rect 201150 2520 201350 2590
rect 201650 2520 201850 2590
rect 202150 2520 202350 2590
rect 202650 2520 202850 2590
rect 203150 2520 203350 2590
rect 203650 2520 203850 2590
rect 204150 2520 204350 2590
rect 204650 2520 204850 2590
rect 205150 2520 205350 2590
rect 205650 2520 205850 2590
rect 206150 2520 206350 2590
rect 206650 2520 206850 2590
rect 207150 2520 207350 2590
rect 207650 2520 207850 2590
rect 198150 2410 198350 2480
rect 198650 2410 198850 2480
rect 199150 2410 199350 2480
rect 199650 2410 199850 2480
rect 200150 2410 200350 2480
rect 200650 2410 200850 2480
rect 201150 2410 201350 2480
rect 201650 2410 201850 2480
rect 202150 2410 202350 2480
rect 202650 2410 202850 2480
rect 203150 2410 203350 2480
rect 203650 2410 203850 2480
rect 204150 2410 204350 2480
rect 204650 2410 204850 2480
rect 205150 2410 205350 2480
rect 205650 2410 205850 2480
rect 206150 2410 206350 2480
rect 206650 2410 206850 2480
rect 207150 2410 207350 2480
rect 207650 2410 207850 2480
rect 198020 2150 198090 2350
rect 198410 2150 198480 2350
rect 198520 2150 198590 2350
rect 198910 2150 198980 2350
rect 199020 2150 199090 2350
rect 199410 2150 199480 2350
rect 199520 2150 199590 2350
rect 199910 2150 199980 2350
rect 200020 2150 200090 2350
rect 200410 2150 200480 2350
rect 200520 2150 200590 2350
rect 200910 2150 200980 2350
rect 201020 2150 201090 2350
rect 201410 2150 201480 2350
rect 201520 2150 201590 2350
rect 201910 2150 201980 2350
rect 202020 2150 202090 2350
rect 202410 2150 202480 2350
rect 202520 2150 202590 2350
rect 202910 2150 202980 2350
rect 203020 2150 203090 2350
rect 203410 2150 203480 2350
rect 203520 2150 203590 2350
rect 203910 2150 203980 2350
rect 204020 2150 204090 2350
rect 204410 2150 204480 2350
rect 204520 2150 204590 2350
rect 204910 2150 204980 2350
rect 205020 2150 205090 2350
rect 205410 2150 205480 2350
rect 205520 2150 205590 2350
rect 205910 2150 205980 2350
rect 206020 2150 206090 2350
rect 206410 2150 206480 2350
rect 206520 2150 206590 2350
rect 206910 2150 206980 2350
rect 207020 2150 207090 2350
rect 207410 2150 207480 2350
rect 207520 2150 207590 2350
rect 207910 2150 207980 2350
rect 198150 2020 198350 2090
rect 198650 2020 198850 2090
rect 199150 2020 199350 2090
rect 199650 2020 199850 2090
rect 200150 2020 200350 2090
rect 200650 2020 200850 2090
rect 201150 2020 201350 2090
rect 201650 2020 201850 2090
rect 202150 2020 202350 2090
rect 202650 2020 202850 2090
rect 203150 2020 203350 2090
rect 203650 2020 203850 2090
rect 204150 2020 204350 2090
rect 204650 2020 204850 2090
rect 205150 2020 205350 2090
rect 205650 2020 205850 2090
rect 206150 2020 206350 2090
rect 206650 2020 206850 2090
rect 207150 2020 207350 2090
rect 207650 2020 207850 2090
<< metal2 >>
rect 250800 136760 251000 136800
rect 250740 136750 251000 136760
rect 250500 135910 250580 135920
rect 250500 135260 250510 135910
rect 250570 135260 250580 135910
rect 250500 135250 250580 135260
rect 250740 134410 250750 136750
rect 250890 134410 251000 136750
rect 250740 134400 251000 134410
rect 171000 121800 182000 122000
rect 171000 119600 171200 121800
rect 181800 119600 182000 121800
rect 171000 119400 182000 119600
rect 222600 121900 232000 122000
rect 222600 119500 222700 121900
rect 231900 119500 232000 121900
rect 222600 119400 232000 119500
rect 181600 119000 182000 119400
rect 231500 119000 232000 119400
rect 196140 103980 196360 104000
rect 196140 103910 196150 103980
rect 196350 103910 196360 103980
rect 196140 103860 196360 103910
rect 196640 103980 196860 104000
rect 196640 103910 196650 103980
rect 196850 103910 196860 103980
rect 196640 103860 196860 103910
rect 197140 103980 197360 104000
rect 197140 103910 197150 103980
rect 197350 103910 197360 103980
rect 197140 103860 197360 103910
rect 197640 103980 197860 104000
rect 197640 103910 197650 103980
rect 197850 103910 197860 103980
rect 197640 103860 197860 103910
rect 198140 103980 198360 104000
rect 198140 103910 198150 103980
rect 198350 103910 198360 103980
rect 198140 103860 198360 103910
rect 198640 103980 198860 104000
rect 198640 103910 198650 103980
rect 198850 103910 198860 103980
rect 198640 103860 198860 103910
rect 199140 103980 199360 104000
rect 199140 103910 199150 103980
rect 199350 103910 199360 103980
rect 199140 103860 199360 103910
rect 199640 103980 199860 104000
rect 199640 103910 199650 103980
rect 199850 103910 199860 103980
rect 199640 103860 199860 103910
rect 200140 103980 200360 104000
rect 200140 103910 200150 103980
rect 200350 103910 200360 103980
rect 200140 103860 200360 103910
rect 200640 103980 200860 104000
rect 200640 103910 200650 103980
rect 200850 103910 200860 103980
rect 200640 103860 200860 103910
rect 201140 103980 201360 104000
rect 201140 103910 201150 103980
rect 201350 103910 201360 103980
rect 201140 103860 201360 103910
rect 201640 103980 201860 104000
rect 201640 103910 201650 103980
rect 201850 103910 201860 103980
rect 201640 103860 201860 103910
rect 202140 103980 202360 104000
rect 202140 103910 202150 103980
rect 202350 103910 202360 103980
rect 202140 103860 202360 103910
rect 202640 103980 202860 104000
rect 202640 103910 202650 103980
rect 202850 103910 202860 103980
rect 202640 103860 202860 103910
rect 203140 103980 203360 104000
rect 203140 103910 203150 103980
rect 203350 103910 203360 103980
rect 203140 103860 203360 103910
rect 203640 103980 203860 104000
rect 203640 103910 203650 103980
rect 203850 103910 203860 103980
rect 203640 103860 203860 103910
rect 204140 103980 204360 104000
rect 204140 103910 204150 103980
rect 204350 103910 204360 103980
rect 204140 103860 204360 103910
rect 204640 103980 204860 104000
rect 204640 103910 204650 103980
rect 204850 103910 204860 103980
rect 204640 103860 204860 103910
rect 205140 103980 205360 104000
rect 205140 103910 205150 103980
rect 205350 103910 205360 103980
rect 205140 103860 205360 103910
rect 205640 103980 205860 104000
rect 205640 103910 205650 103980
rect 205850 103910 205860 103980
rect 205640 103860 205860 103910
rect 206140 103980 206360 104000
rect 206140 103910 206150 103980
rect 206350 103910 206360 103980
rect 206140 103860 206360 103910
rect 206640 103980 206860 104000
rect 206640 103910 206650 103980
rect 206850 103910 206860 103980
rect 206640 103860 206860 103910
rect 207140 103980 207360 104000
rect 207140 103910 207150 103980
rect 207350 103910 207360 103980
rect 207140 103860 207360 103910
rect 207640 103980 207860 104000
rect 207640 103910 207650 103980
rect 207850 103910 207860 103980
rect 207640 103860 207860 103910
rect 196000 103850 208000 103860
rect 196000 103650 196020 103850
rect 196090 103650 196410 103850
rect 196480 103650 196520 103850
rect 196590 103650 196910 103850
rect 196980 103650 197020 103850
rect 197090 103650 197410 103850
rect 197480 103650 197520 103850
rect 197590 103650 197910 103850
rect 197980 103650 198020 103850
rect 198090 103650 198410 103850
rect 198480 103650 198520 103850
rect 198590 103650 198910 103850
rect 198980 103650 199020 103850
rect 199090 103650 199410 103850
rect 199480 103650 199520 103850
rect 199590 103650 199910 103850
rect 199980 103650 200020 103850
rect 200090 103650 200410 103850
rect 200480 103650 200520 103850
rect 200590 103650 200910 103850
rect 200980 103650 201020 103850
rect 201090 103650 201410 103850
rect 201480 103650 201520 103850
rect 201590 103650 201910 103850
rect 201980 103650 202020 103850
rect 202090 103650 202410 103850
rect 202480 103650 202520 103850
rect 202590 103650 202910 103850
rect 202980 103650 203020 103850
rect 203090 103650 203410 103850
rect 203480 103650 203520 103850
rect 203590 103650 203910 103850
rect 203980 103650 204020 103850
rect 204090 103650 204410 103850
rect 204480 103650 204520 103850
rect 204590 103650 204910 103850
rect 204980 103650 205020 103850
rect 205090 103650 205410 103850
rect 205480 103650 205520 103850
rect 205590 103650 205910 103850
rect 205980 103650 206020 103850
rect 206090 103650 206410 103850
rect 206480 103650 206520 103850
rect 206590 103650 206910 103850
rect 206980 103650 207020 103850
rect 207090 103650 207410 103850
rect 207480 103650 207520 103850
rect 207590 103650 207910 103850
rect 207980 103650 208000 103850
rect 196000 103640 208000 103650
rect 196140 103590 196360 103640
rect 196140 103520 196150 103590
rect 196350 103520 196360 103590
rect 196140 103480 196360 103520
rect 196140 103410 196150 103480
rect 196350 103410 196360 103480
rect 196140 103360 196360 103410
rect 196640 103590 196860 103640
rect 196640 103520 196650 103590
rect 196850 103520 196860 103590
rect 196640 103480 196860 103520
rect 196640 103410 196650 103480
rect 196850 103410 196860 103480
rect 196640 103360 196860 103410
rect 197140 103590 197360 103640
rect 197140 103520 197150 103590
rect 197350 103520 197360 103590
rect 197140 103480 197360 103520
rect 197140 103410 197150 103480
rect 197350 103410 197360 103480
rect 197140 103360 197360 103410
rect 197640 103590 197860 103640
rect 197640 103520 197650 103590
rect 197850 103520 197860 103590
rect 197640 103480 197860 103520
rect 197640 103410 197650 103480
rect 197850 103410 197860 103480
rect 197640 103360 197860 103410
rect 198140 103590 198360 103640
rect 198140 103520 198150 103590
rect 198350 103520 198360 103590
rect 198140 103480 198360 103520
rect 198140 103410 198150 103480
rect 198350 103410 198360 103480
rect 198140 103360 198360 103410
rect 198640 103590 198860 103640
rect 198640 103520 198650 103590
rect 198850 103520 198860 103590
rect 198640 103480 198860 103520
rect 198640 103410 198650 103480
rect 198850 103410 198860 103480
rect 198640 103360 198860 103410
rect 199140 103590 199360 103640
rect 199140 103520 199150 103590
rect 199350 103520 199360 103590
rect 199140 103480 199360 103520
rect 199140 103410 199150 103480
rect 199350 103410 199360 103480
rect 199140 103360 199360 103410
rect 199640 103590 199860 103640
rect 199640 103520 199650 103590
rect 199850 103520 199860 103590
rect 199640 103480 199860 103520
rect 199640 103410 199650 103480
rect 199850 103410 199860 103480
rect 199640 103360 199860 103410
rect 200140 103590 200360 103640
rect 200140 103520 200150 103590
rect 200350 103520 200360 103590
rect 200140 103480 200360 103520
rect 200140 103410 200150 103480
rect 200350 103410 200360 103480
rect 200140 103360 200360 103410
rect 200640 103590 200860 103640
rect 200640 103520 200650 103590
rect 200850 103520 200860 103590
rect 200640 103480 200860 103520
rect 200640 103410 200650 103480
rect 200850 103410 200860 103480
rect 200640 103360 200860 103410
rect 201140 103590 201360 103640
rect 201140 103520 201150 103590
rect 201350 103520 201360 103590
rect 201140 103480 201360 103520
rect 201140 103410 201150 103480
rect 201350 103410 201360 103480
rect 201140 103360 201360 103410
rect 201640 103590 201860 103640
rect 201640 103520 201650 103590
rect 201850 103520 201860 103590
rect 201640 103480 201860 103520
rect 201640 103410 201650 103480
rect 201850 103410 201860 103480
rect 201640 103360 201860 103410
rect 202140 103590 202360 103640
rect 202140 103520 202150 103590
rect 202350 103520 202360 103590
rect 202140 103480 202360 103520
rect 202140 103410 202150 103480
rect 202350 103410 202360 103480
rect 202140 103360 202360 103410
rect 202640 103590 202860 103640
rect 202640 103520 202650 103590
rect 202850 103520 202860 103590
rect 202640 103480 202860 103520
rect 202640 103410 202650 103480
rect 202850 103410 202860 103480
rect 202640 103360 202860 103410
rect 203140 103590 203360 103640
rect 203140 103520 203150 103590
rect 203350 103520 203360 103590
rect 203140 103480 203360 103520
rect 203140 103410 203150 103480
rect 203350 103410 203360 103480
rect 203140 103360 203360 103410
rect 203640 103590 203860 103640
rect 203640 103520 203650 103590
rect 203850 103520 203860 103590
rect 203640 103480 203860 103520
rect 203640 103410 203650 103480
rect 203850 103410 203860 103480
rect 203640 103360 203860 103410
rect 204140 103590 204360 103640
rect 204140 103520 204150 103590
rect 204350 103520 204360 103590
rect 204140 103480 204360 103520
rect 204140 103410 204150 103480
rect 204350 103410 204360 103480
rect 204140 103360 204360 103410
rect 204640 103590 204860 103640
rect 204640 103520 204650 103590
rect 204850 103520 204860 103590
rect 204640 103480 204860 103520
rect 204640 103410 204650 103480
rect 204850 103410 204860 103480
rect 204640 103360 204860 103410
rect 205140 103590 205360 103640
rect 205140 103520 205150 103590
rect 205350 103520 205360 103590
rect 205140 103480 205360 103520
rect 205140 103410 205150 103480
rect 205350 103410 205360 103480
rect 205140 103360 205360 103410
rect 205640 103590 205860 103640
rect 205640 103520 205650 103590
rect 205850 103520 205860 103590
rect 205640 103480 205860 103520
rect 205640 103410 205650 103480
rect 205850 103410 205860 103480
rect 205640 103360 205860 103410
rect 206140 103590 206360 103640
rect 206140 103520 206150 103590
rect 206350 103520 206360 103590
rect 206140 103480 206360 103520
rect 206140 103410 206150 103480
rect 206350 103410 206360 103480
rect 206140 103360 206360 103410
rect 206640 103590 206860 103640
rect 206640 103520 206650 103590
rect 206850 103520 206860 103590
rect 206640 103480 206860 103520
rect 206640 103410 206650 103480
rect 206850 103410 206860 103480
rect 206640 103360 206860 103410
rect 207140 103590 207360 103640
rect 207140 103520 207150 103590
rect 207350 103520 207360 103590
rect 207140 103480 207360 103520
rect 207140 103410 207150 103480
rect 207350 103410 207360 103480
rect 207140 103360 207360 103410
rect 207640 103590 207860 103640
rect 207640 103520 207650 103590
rect 207850 103520 207860 103590
rect 207640 103480 207860 103520
rect 207640 103410 207650 103480
rect 207850 103410 207860 103480
rect 207640 103360 207860 103410
rect 196000 103350 208000 103360
rect 196000 103150 196020 103350
rect 196090 103150 196410 103350
rect 196480 103150 196520 103350
rect 196590 103150 196910 103350
rect 196980 103150 197020 103350
rect 197090 103150 197410 103350
rect 197480 103150 197520 103350
rect 197590 103150 197910 103350
rect 197980 103150 198020 103350
rect 198090 103150 198410 103350
rect 198480 103150 198520 103350
rect 198590 103150 198910 103350
rect 198980 103150 199020 103350
rect 199090 103150 199410 103350
rect 199480 103150 199520 103350
rect 199590 103150 199910 103350
rect 199980 103150 200020 103350
rect 200090 103150 200410 103350
rect 200480 103150 200520 103350
rect 200590 103150 200910 103350
rect 200980 103150 201020 103350
rect 201090 103150 201410 103350
rect 201480 103150 201520 103350
rect 201590 103150 201910 103350
rect 201980 103150 202020 103350
rect 202090 103150 202410 103350
rect 202480 103150 202520 103350
rect 202590 103150 202910 103350
rect 202980 103150 203020 103350
rect 203090 103150 203410 103350
rect 203480 103150 203520 103350
rect 203590 103150 203910 103350
rect 203980 103150 204020 103350
rect 204090 103150 204410 103350
rect 204480 103150 204520 103350
rect 204590 103150 204910 103350
rect 204980 103150 205020 103350
rect 205090 103150 205410 103350
rect 205480 103150 205520 103350
rect 205590 103150 205910 103350
rect 205980 103150 206020 103350
rect 206090 103150 206410 103350
rect 206480 103150 206520 103350
rect 206590 103150 206910 103350
rect 206980 103150 207020 103350
rect 207090 103150 207410 103350
rect 207480 103150 207520 103350
rect 207590 103150 207910 103350
rect 207980 103150 208000 103350
rect 196000 103140 208000 103150
rect 196140 103090 196360 103140
rect 196140 103020 196150 103090
rect 196350 103020 196360 103090
rect 196140 102980 196360 103020
rect 196140 102910 196150 102980
rect 196350 102910 196360 102980
rect 196140 102860 196360 102910
rect 196640 103090 196860 103140
rect 196640 103020 196650 103090
rect 196850 103020 196860 103090
rect 196640 102980 196860 103020
rect 196640 102910 196650 102980
rect 196850 102910 196860 102980
rect 196640 102860 196860 102910
rect 197140 103090 197360 103140
rect 197140 103020 197150 103090
rect 197350 103020 197360 103090
rect 197140 102980 197360 103020
rect 197140 102910 197150 102980
rect 197350 102910 197360 102980
rect 197140 102860 197360 102910
rect 197640 103090 197860 103140
rect 197640 103020 197650 103090
rect 197850 103020 197860 103090
rect 197640 102980 197860 103020
rect 197640 102910 197650 102980
rect 197850 102910 197860 102980
rect 197640 102860 197860 102910
rect 198140 103090 198360 103140
rect 198140 103020 198150 103090
rect 198350 103020 198360 103090
rect 198140 102980 198360 103020
rect 198140 102910 198150 102980
rect 198350 102910 198360 102980
rect 198140 102860 198360 102910
rect 198640 103090 198860 103140
rect 198640 103020 198650 103090
rect 198850 103020 198860 103090
rect 198640 102980 198860 103020
rect 198640 102910 198650 102980
rect 198850 102910 198860 102980
rect 198640 102860 198860 102910
rect 199140 103090 199360 103140
rect 199140 103020 199150 103090
rect 199350 103020 199360 103090
rect 199140 102980 199360 103020
rect 199140 102910 199150 102980
rect 199350 102910 199360 102980
rect 199140 102860 199360 102910
rect 199640 103090 199860 103140
rect 199640 103020 199650 103090
rect 199850 103020 199860 103090
rect 199640 102980 199860 103020
rect 199640 102910 199650 102980
rect 199850 102910 199860 102980
rect 199640 102860 199860 102910
rect 200140 103090 200360 103140
rect 200140 103020 200150 103090
rect 200350 103020 200360 103090
rect 200140 102980 200360 103020
rect 200140 102910 200150 102980
rect 200350 102910 200360 102980
rect 200140 102860 200360 102910
rect 200640 103090 200860 103140
rect 200640 103020 200650 103090
rect 200850 103020 200860 103090
rect 200640 102980 200860 103020
rect 200640 102910 200650 102980
rect 200850 102910 200860 102980
rect 200640 102860 200860 102910
rect 201140 103090 201360 103140
rect 201140 103020 201150 103090
rect 201350 103020 201360 103090
rect 201140 102980 201360 103020
rect 201140 102910 201150 102980
rect 201350 102910 201360 102980
rect 201140 102860 201360 102910
rect 201640 103090 201860 103140
rect 201640 103020 201650 103090
rect 201850 103020 201860 103090
rect 201640 102980 201860 103020
rect 201640 102910 201650 102980
rect 201850 102910 201860 102980
rect 201640 102860 201860 102910
rect 202140 103090 202360 103140
rect 202140 103020 202150 103090
rect 202350 103020 202360 103090
rect 202140 102980 202360 103020
rect 202140 102910 202150 102980
rect 202350 102910 202360 102980
rect 202140 102860 202360 102910
rect 202640 103090 202860 103140
rect 202640 103020 202650 103090
rect 202850 103020 202860 103090
rect 202640 102980 202860 103020
rect 202640 102910 202650 102980
rect 202850 102910 202860 102980
rect 202640 102860 202860 102910
rect 203140 103090 203360 103140
rect 203140 103020 203150 103090
rect 203350 103020 203360 103090
rect 203140 102980 203360 103020
rect 203140 102910 203150 102980
rect 203350 102910 203360 102980
rect 203140 102860 203360 102910
rect 203640 103090 203860 103140
rect 203640 103020 203650 103090
rect 203850 103020 203860 103090
rect 203640 102980 203860 103020
rect 203640 102910 203650 102980
rect 203850 102910 203860 102980
rect 203640 102860 203860 102910
rect 204140 103090 204360 103140
rect 204140 103020 204150 103090
rect 204350 103020 204360 103090
rect 204140 102980 204360 103020
rect 204140 102910 204150 102980
rect 204350 102910 204360 102980
rect 204140 102860 204360 102910
rect 204640 103090 204860 103140
rect 204640 103020 204650 103090
rect 204850 103020 204860 103090
rect 204640 102980 204860 103020
rect 204640 102910 204650 102980
rect 204850 102910 204860 102980
rect 204640 102860 204860 102910
rect 205140 103090 205360 103140
rect 205140 103020 205150 103090
rect 205350 103020 205360 103090
rect 205140 102980 205360 103020
rect 205140 102910 205150 102980
rect 205350 102910 205360 102980
rect 205140 102860 205360 102910
rect 205640 103090 205860 103140
rect 205640 103020 205650 103090
rect 205850 103020 205860 103090
rect 205640 102980 205860 103020
rect 205640 102910 205650 102980
rect 205850 102910 205860 102980
rect 205640 102860 205860 102910
rect 206140 103090 206360 103140
rect 206140 103020 206150 103090
rect 206350 103020 206360 103090
rect 206140 102980 206360 103020
rect 206140 102910 206150 102980
rect 206350 102910 206360 102980
rect 206140 102860 206360 102910
rect 206640 103090 206860 103140
rect 206640 103020 206650 103090
rect 206850 103020 206860 103090
rect 206640 102980 206860 103020
rect 206640 102910 206650 102980
rect 206850 102910 206860 102980
rect 206640 102860 206860 102910
rect 207140 103090 207360 103140
rect 207140 103020 207150 103090
rect 207350 103020 207360 103090
rect 207140 102980 207360 103020
rect 207140 102910 207150 102980
rect 207350 102910 207360 102980
rect 207140 102860 207360 102910
rect 207640 103090 207860 103140
rect 207640 103020 207650 103090
rect 207850 103020 207860 103090
rect 207640 102980 207860 103020
rect 207640 102910 207650 102980
rect 207850 102910 207860 102980
rect 207640 102860 207860 102910
rect 196000 102850 208000 102860
rect 196000 102650 196020 102850
rect 196090 102650 196410 102850
rect 196480 102650 196520 102850
rect 196590 102650 196910 102850
rect 196980 102650 197020 102850
rect 197090 102650 197410 102850
rect 197480 102650 197520 102850
rect 197590 102650 197910 102850
rect 197980 102650 198020 102850
rect 198090 102650 198410 102850
rect 198480 102650 198520 102850
rect 198590 102650 198910 102850
rect 198980 102650 199020 102850
rect 199090 102650 199410 102850
rect 199480 102650 199520 102850
rect 199590 102650 199910 102850
rect 199980 102650 200020 102850
rect 200090 102650 200410 102850
rect 200480 102650 200520 102850
rect 200590 102650 200910 102850
rect 200980 102650 201020 102850
rect 201090 102650 201410 102850
rect 201480 102650 201520 102850
rect 201590 102650 201910 102850
rect 201980 102650 202020 102850
rect 202090 102650 202410 102850
rect 202480 102650 202520 102850
rect 202590 102650 202910 102850
rect 202980 102650 203020 102850
rect 203090 102650 203410 102850
rect 203480 102650 203520 102850
rect 203590 102650 203910 102850
rect 203980 102650 204020 102850
rect 204090 102650 204410 102850
rect 204480 102650 204520 102850
rect 204590 102650 204910 102850
rect 204980 102650 205020 102850
rect 205090 102650 205410 102850
rect 205480 102650 205520 102850
rect 205590 102650 205910 102850
rect 205980 102650 206020 102850
rect 206090 102650 206410 102850
rect 206480 102650 206520 102850
rect 206590 102650 206910 102850
rect 206980 102650 207020 102850
rect 207090 102650 207410 102850
rect 207480 102650 207520 102850
rect 207590 102650 207910 102850
rect 207980 102650 208000 102850
rect 196000 102640 208000 102650
rect 196140 102590 196360 102640
rect 196140 102520 196150 102590
rect 196350 102520 196360 102590
rect 196140 102480 196360 102520
rect 196140 102410 196150 102480
rect 196350 102410 196360 102480
rect 196140 102360 196360 102410
rect 196640 102590 196860 102640
rect 196640 102520 196650 102590
rect 196850 102520 196860 102590
rect 196640 102480 196860 102520
rect 196640 102410 196650 102480
rect 196850 102410 196860 102480
rect 196640 102360 196860 102410
rect 197140 102590 197360 102640
rect 197140 102520 197150 102590
rect 197350 102520 197360 102590
rect 197140 102480 197360 102520
rect 197140 102410 197150 102480
rect 197350 102410 197360 102480
rect 197140 102360 197360 102410
rect 197640 102590 197860 102640
rect 197640 102520 197650 102590
rect 197850 102520 197860 102590
rect 197640 102480 197860 102520
rect 197640 102410 197650 102480
rect 197850 102410 197860 102480
rect 197640 102360 197860 102410
rect 198140 102590 198360 102640
rect 198140 102520 198150 102590
rect 198350 102520 198360 102590
rect 198140 102480 198360 102520
rect 198140 102410 198150 102480
rect 198350 102410 198360 102480
rect 198140 102360 198360 102410
rect 198640 102590 198860 102640
rect 198640 102520 198650 102590
rect 198850 102520 198860 102590
rect 198640 102480 198860 102520
rect 198640 102410 198650 102480
rect 198850 102410 198860 102480
rect 198640 102360 198860 102410
rect 199140 102590 199360 102640
rect 199140 102520 199150 102590
rect 199350 102520 199360 102590
rect 199140 102480 199360 102520
rect 199140 102410 199150 102480
rect 199350 102410 199360 102480
rect 199140 102360 199360 102410
rect 199640 102590 199860 102640
rect 199640 102520 199650 102590
rect 199850 102520 199860 102590
rect 199640 102480 199860 102520
rect 199640 102410 199650 102480
rect 199850 102410 199860 102480
rect 199640 102360 199860 102410
rect 200140 102590 200360 102640
rect 200140 102520 200150 102590
rect 200350 102520 200360 102590
rect 200140 102480 200360 102520
rect 200140 102410 200150 102480
rect 200350 102410 200360 102480
rect 200140 102360 200360 102410
rect 200640 102590 200860 102640
rect 200640 102520 200650 102590
rect 200850 102520 200860 102590
rect 200640 102480 200860 102520
rect 200640 102410 200650 102480
rect 200850 102410 200860 102480
rect 200640 102360 200860 102410
rect 201140 102590 201360 102640
rect 201140 102520 201150 102590
rect 201350 102520 201360 102590
rect 201140 102480 201360 102520
rect 201140 102410 201150 102480
rect 201350 102410 201360 102480
rect 201140 102360 201360 102410
rect 201640 102590 201860 102640
rect 201640 102520 201650 102590
rect 201850 102520 201860 102590
rect 201640 102480 201860 102520
rect 201640 102410 201650 102480
rect 201850 102410 201860 102480
rect 201640 102360 201860 102410
rect 202140 102590 202360 102640
rect 202140 102520 202150 102590
rect 202350 102520 202360 102590
rect 202140 102480 202360 102520
rect 202140 102410 202150 102480
rect 202350 102410 202360 102480
rect 202140 102360 202360 102410
rect 202640 102590 202860 102640
rect 202640 102520 202650 102590
rect 202850 102520 202860 102590
rect 202640 102480 202860 102520
rect 202640 102410 202650 102480
rect 202850 102410 202860 102480
rect 202640 102360 202860 102410
rect 203140 102590 203360 102640
rect 203140 102520 203150 102590
rect 203350 102520 203360 102590
rect 203140 102480 203360 102520
rect 203140 102410 203150 102480
rect 203350 102410 203360 102480
rect 203140 102360 203360 102410
rect 203640 102590 203860 102640
rect 203640 102520 203650 102590
rect 203850 102520 203860 102590
rect 203640 102480 203860 102520
rect 203640 102410 203650 102480
rect 203850 102410 203860 102480
rect 203640 102360 203860 102410
rect 204140 102590 204360 102640
rect 204140 102520 204150 102590
rect 204350 102520 204360 102590
rect 204140 102480 204360 102520
rect 204140 102410 204150 102480
rect 204350 102410 204360 102480
rect 204140 102360 204360 102410
rect 204640 102590 204860 102640
rect 204640 102520 204650 102590
rect 204850 102520 204860 102590
rect 204640 102480 204860 102520
rect 204640 102410 204650 102480
rect 204850 102410 204860 102480
rect 204640 102360 204860 102410
rect 205140 102590 205360 102640
rect 205140 102520 205150 102590
rect 205350 102520 205360 102590
rect 205140 102480 205360 102520
rect 205140 102410 205150 102480
rect 205350 102410 205360 102480
rect 205140 102360 205360 102410
rect 205640 102590 205860 102640
rect 205640 102520 205650 102590
rect 205850 102520 205860 102590
rect 205640 102480 205860 102520
rect 205640 102410 205650 102480
rect 205850 102410 205860 102480
rect 205640 102360 205860 102410
rect 206140 102590 206360 102640
rect 206140 102520 206150 102590
rect 206350 102520 206360 102590
rect 206140 102480 206360 102520
rect 206140 102410 206150 102480
rect 206350 102410 206360 102480
rect 206140 102360 206360 102410
rect 206640 102590 206860 102640
rect 206640 102520 206650 102590
rect 206850 102520 206860 102590
rect 206640 102480 206860 102520
rect 206640 102410 206650 102480
rect 206850 102410 206860 102480
rect 206640 102360 206860 102410
rect 207140 102590 207360 102640
rect 207140 102520 207150 102590
rect 207350 102520 207360 102590
rect 207140 102480 207360 102520
rect 207140 102410 207150 102480
rect 207350 102410 207360 102480
rect 207140 102360 207360 102410
rect 207640 102590 207860 102640
rect 207640 102520 207650 102590
rect 207850 102520 207860 102590
rect 207640 102480 207860 102520
rect 207640 102410 207650 102480
rect 207850 102410 207860 102480
rect 207640 102360 207860 102410
rect 196000 102350 208000 102360
rect 196000 102150 196020 102350
rect 196090 102150 196410 102350
rect 196480 102150 196520 102350
rect 196590 102150 196910 102350
rect 196980 102150 197020 102350
rect 197090 102150 197410 102350
rect 197480 102150 197520 102350
rect 197590 102150 197910 102350
rect 197980 102150 198020 102350
rect 198090 102150 198410 102350
rect 198480 102150 198520 102350
rect 198590 102150 198910 102350
rect 198980 102150 199020 102350
rect 199090 102150 199410 102350
rect 199480 102150 199520 102350
rect 199590 102150 199910 102350
rect 199980 102150 200020 102350
rect 200090 102150 200410 102350
rect 200480 102150 200520 102350
rect 200590 102150 200910 102350
rect 200980 102150 201020 102350
rect 201090 102150 201410 102350
rect 201480 102150 201520 102350
rect 201590 102150 201910 102350
rect 201980 102150 202020 102350
rect 202090 102150 202410 102350
rect 202480 102150 202520 102350
rect 202590 102150 202910 102350
rect 202980 102150 203020 102350
rect 203090 102150 203410 102350
rect 203480 102150 203520 102350
rect 203590 102150 203910 102350
rect 203980 102150 204020 102350
rect 204090 102150 204410 102350
rect 204480 102150 204520 102350
rect 204590 102150 204910 102350
rect 204980 102150 205020 102350
rect 205090 102150 205410 102350
rect 205480 102150 205520 102350
rect 205590 102150 205910 102350
rect 205980 102150 206020 102350
rect 206090 102150 206410 102350
rect 206480 102150 206520 102350
rect 206590 102150 206910 102350
rect 206980 102150 207020 102350
rect 207090 102150 207410 102350
rect 207480 102150 207520 102350
rect 207590 102150 207910 102350
rect 207980 102150 208000 102350
rect 196000 102140 208000 102150
rect 196140 102090 196360 102140
rect 196140 102020 196150 102090
rect 196350 102020 196360 102090
rect 196140 101980 196360 102020
rect 196140 101910 196150 101980
rect 196350 101910 196360 101980
rect 196140 101860 196360 101910
rect 196640 102090 196860 102140
rect 196640 102020 196650 102090
rect 196850 102020 196860 102090
rect 196640 101980 196860 102020
rect 196640 101910 196650 101980
rect 196850 101910 196860 101980
rect 196640 101860 196860 101910
rect 197140 102090 197360 102140
rect 197140 102020 197150 102090
rect 197350 102020 197360 102090
rect 197140 101980 197360 102020
rect 197140 101910 197150 101980
rect 197350 101910 197360 101980
rect 197140 101860 197360 101910
rect 197640 102090 197860 102140
rect 197640 102020 197650 102090
rect 197850 102020 197860 102090
rect 197640 101980 197860 102020
rect 197640 101910 197650 101980
rect 197850 101910 197860 101980
rect 197640 101860 197860 101910
rect 198140 102090 198360 102140
rect 198140 102020 198150 102090
rect 198350 102020 198360 102090
rect 198140 101980 198360 102020
rect 198140 101910 198150 101980
rect 198350 101910 198360 101980
rect 198140 101860 198360 101910
rect 198640 102090 198860 102140
rect 198640 102020 198650 102090
rect 198850 102020 198860 102090
rect 198640 101980 198860 102020
rect 198640 101910 198650 101980
rect 198850 101910 198860 101980
rect 198640 101860 198860 101910
rect 199140 102090 199360 102140
rect 199140 102020 199150 102090
rect 199350 102020 199360 102090
rect 199140 101980 199360 102020
rect 199140 101910 199150 101980
rect 199350 101910 199360 101980
rect 199140 101860 199360 101910
rect 199640 102090 199860 102140
rect 199640 102020 199650 102090
rect 199850 102020 199860 102090
rect 199640 101980 199860 102020
rect 199640 101910 199650 101980
rect 199850 101910 199860 101980
rect 199640 101860 199860 101910
rect 200140 102090 200360 102140
rect 200140 102020 200150 102090
rect 200350 102020 200360 102090
rect 200140 101980 200360 102020
rect 200140 101910 200150 101980
rect 200350 101910 200360 101980
rect 200140 101860 200360 101910
rect 200640 102090 200860 102140
rect 200640 102020 200650 102090
rect 200850 102020 200860 102090
rect 200640 101980 200860 102020
rect 200640 101910 200650 101980
rect 200850 101910 200860 101980
rect 200640 101860 200860 101910
rect 201140 102090 201360 102140
rect 201140 102020 201150 102090
rect 201350 102020 201360 102090
rect 201140 101980 201360 102020
rect 201140 101910 201150 101980
rect 201350 101910 201360 101980
rect 201140 101860 201360 101910
rect 201640 102090 201860 102140
rect 201640 102020 201650 102090
rect 201850 102020 201860 102090
rect 201640 101980 201860 102020
rect 201640 101910 201650 101980
rect 201850 101910 201860 101980
rect 201640 101860 201860 101910
rect 202140 102090 202360 102140
rect 202140 102020 202150 102090
rect 202350 102020 202360 102090
rect 202140 101980 202360 102020
rect 202140 101910 202150 101980
rect 202350 101910 202360 101980
rect 202140 101860 202360 101910
rect 202640 102090 202860 102140
rect 202640 102020 202650 102090
rect 202850 102020 202860 102090
rect 202640 101980 202860 102020
rect 202640 101910 202650 101980
rect 202850 101910 202860 101980
rect 202640 101860 202860 101910
rect 203140 102090 203360 102140
rect 203140 102020 203150 102090
rect 203350 102020 203360 102090
rect 203140 101980 203360 102020
rect 203140 101910 203150 101980
rect 203350 101910 203360 101980
rect 203140 101860 203360 101910
rect 203640 102090 203860 102140
rect 203640 102020 203650 102090
rect 203850 102020 203860 102090
rect 203640 101980 203860 102020
rect 203640 101910 203650 101980
rect 203850 101910 203860 101980
rect 203640 101860 203860 101910
rect 204140 102090 204360 102140
rect 204140 102020 204150 102090
rect 204350 102020 204360 102090
rect 204140 101980 204360 102020
rect 204140 101910 204150 101980
rect 204350 101910 204360 101980
rect 204140 101860 204360 101910
rect 204640 102090 204860 102140
rect 204640 102020 204650 102090
rect 204850 102020 204860 102090
rect 204640 101980 204860 102020
rect 204640 101910 204650 101980
rect 204850 101910 204860 101980
rect 204640 101860 204860 101910
rect 205140 102090 205360 102140
rect 205140 102020 205150 102090
rect 205350 102020 205360 102090
rect 205140 101980 205360 102020
rect 205140 101910 205150 101980
rect 205350 101910 205360 101980
rect 205140 101860 205360 101910
rect 205640 102090 205860 102140
rect 205640 102020 205650 102090
rect 205850 102020 205860 102090
rect 205640 101980 205860 102020
rect 205640 101910 205650 101980
rect 205850 101910 205860 101980
rect 205640 101860 205860 101910
rect 206140 102090 206360 102140
rect 206140 102020 206150 102090
rect 206350 102020 206360 102090
rect 206140 101980 206360 102020
rect 206140 101910 206150 101980
rect 206350 101910 206360 101980
rect 206140 101860 206360 101910
rect 206640 102090 206860 102140
rect 206640 102020 206650 102090
rect 206850 102020 206860 102090
rect 206640 101980 206860 102020
rect 206640 101910 206650 101980
rect 206850 101910 206860 101980
rect 206640 101860 206860 101910
rect 207140 102090 207360 102140
rect 207140 102020 207150 102090
rect 207350 102020 207360 102090
rect 207140 101980 207360 102020
rect 207140 101910 207150 101980
rect 207350 101910 207360 101980
rect 207140 101860 207360 101910
rect 207640 102090 207860 102140
rect 207640 102020 207650 102090
rect 207850 102020 207860 102090
rect 207640 101980 207860 102020
rect 207640 101910 207650 101980
rect 207850 101910 207860 101980
rect 207640 101860 207860 101910
rect 196000 101850 208000 101860
rect 196000 101650 196020 101850
rect 196090 101650 196410 101850
rect 196480 101650 196520 101850
rect 196590 101650 196910 101850
rect 196980 101650 197020 101850
rect 197090 101650 197410 101850
rect 197480 101650 197520 101850
rect 197590 101650 197910 101850
rect 197980 101650 198020 101850
rect 198090 101650 198410 101850
rect 198480 101650 198520 101850
rect 198590 101650 198910 101850
rect 198980 101650 199020 101850
rect 199090 101650 199410 101850
rect 199480 101650 199520 101850
rect 199590 101650 199910 101850
rect 199980 101650 200020 101850
rect 200090 101650 200410 101850
rect 200480 101650 200520 101850
rect 200590 101650 200910 101850
rect 200980 101650 201020 101850
rect 201090 101650 201410 101850
rect 201480 101650 201520 101850
rect 201590 101650 201910 101850
rect 201980 101650 202020 101850
rect 202090 101650 202410 101850
rect 202480 101650 202520 101850
rect 202590 101650 202910 101850
rect 202980 101650 203020 101850
rect 203090 101650 203410 101850
rect 203480 101650 203520 101850
rect 203590 101650 203910 101850
rect 203980 101650 204020 101850
rect 204090 101650 204410 101850
rect 204480 101650 204520 101850
rect 204590 101650 204910 101850
rect 204980 101650 205020 101850
rect 205090 101650 205410 101850
rect 205480 101650 205520 101850
rect 205590 101650 205910 101850
rect 205980 101650 206020 101850
rect 206090 101650 206410 101850
rect 206480 101650 206520 101850
rect 206590 101650 206910 101850
rect 206980 101650 207020 101850
rect 207090 101650 207410 101850
rect 207480 101650 207520 101850
rect 207590 101650 207910 101850
rect 207980 101650 208000 101850
rect 196000 101640 208000 101650
rect 196140 101590 196360 101640
rect 196140 101520 196150 101590
rect 196350 101520 196360 101590
rect 196140 101480 196360 101520
rect 196140 101410 196150 101480
rect 196350 101410 196360 101480
rect 196140 101360 196360 101410
rect 196640 101590 196860 101640
rect 196640 101520 196650 101590
rect 196850 101520 196860 101590
rect 196640 101480 196860 101520
rect 196640 101410 196650 101480
rect 196850 101410 196860 101480
rect 196640 101360 196860 101410
rect 197140 101590 197360 101640
rect 197140 101520 197150 101590
rect 197350 101520 197360 101590
rect 197140 101480 197360 101520
rect 197140 101410 197150 101480
rect 197350 101410 197360 101480
rect 197140 101360 197360 101410
rect 197640 101590 197860 101640
rect 197640 101520 197650 101590
rect 197850 101520 197860 101590
rect 197640 101480 197860 101520
rect 197640 101410 197650 101480
rect 197850 101410 197860 101480
rect 197640 101360 197860 101410
rect 198140 101590 198360 101640
rect 198140 101520 198150 101590
rect 198350 101520 198360 101590
rect 198140 101480 198360 101520
rect 198140 101410 198150 101480
rect 198350 101410 198360 101480
rect 198140 101360 198360 101410
rect 198640 101590 198860 101640
rect 198640 101520 198650 101590
rect 198850 101520 198860 101590
rect 198640 101480 198860 101520
rect 198640 101410 198650 101480
rect 198850 101410 198860 101480
rect 198640 101360 198860 101410
rect 199140 101590 199360 101640
rect 199140 101520 199150 101590
rect 199350 101520 199360 101590
rect 199140 101480 199360 101520
rect 199140 101410 199150 101480
rect 199350 101410 199360 101480
rect 199140 101360 199360 101410
rect 199640 101590 199860 101640
rect 199640 101520 199650 101590
rect 199850 101520 199860 101590
rect 199640 101480 199860 101520
rect 199640 101410 199650 101480
rect 199850 101410 199860 101480
rect 199640 101360 199860 101410
rect 200140 101590 200360 101640
rect 200140 101520 200150 101590
rect 200350 101520 200360 101590
rect 200140 101480 200360 101520
rect 200140 101410 200150 101480
rect 200350 101410 200360 101480
rect 200140 101360 200360 101410
rect 200640 101590 200860 101640
rect 200640 101520 200650 101590
rect 200850 101520 200860 101590
rect 200640 101480 200860 101520
rect 200640 101410 200650 101480
rect 200850 101410 200860 101480
rect 200640 101360 200860 101410
rect 201140 101590 201360 101640
rect 201140 101520 201150 101590
rect 201350 101520 201360 101590
rect 201140 101480 201360 101520
rect 201140 101410 201150 101480
rect 201350 101410 201360 101480
rect 201140 101360 201360 101410
rect 201640 101590 201860 101640
rect 201640 101520 201650 101590
rect 201850 101520 201860 101590
rect 201640 101480 201860 101520
rect 201640 101410 201650 101480
rect 201850 101410 201860 101480
rect 201640 101360 201860 101410
rect 202140 101590 202360 101640
rect 202140 101520 202150 101590
rect 202350 101520 202360 101590
rect 202140 101480 202360 101520
rect 202140 101410 202150 101480
rect 202350 101410 202360 101480
rect 202140 101360 202360 101410
rect 202640 101590 202860 101640
rect 202640 101520 202650 101590
rect 202850 101520 202860 101590
rect 202640 101480 202860 101520
rect 202640 101410 202650 101480
rect 202850 101410 202860 101480
rect 202640 101360 202860 101410
rect 203140 101590 203360 101640
rect 203140 101520 203150 101590
rect 203350 101520 203360 101590
rect 203140 101480 203360 101520
rect 203140 101410 203150 101480
rect 203350 101410 203360 101480
rect 203140 101360 203360 101410
rect 203640 101590 203860 101640
rect 203640 101520 203650 101590
rect 203850 101520 203860 101590
rect 203640 101480 203860 101520
rect 203640 101410 203650 101480
rect 203850 101410 203860 101480
rect 203640 101360 203860 101410
rect 204140 101590 204360 101640
rect 204140 101520 204150 101590
rect 204350 101520 204360 101590
rect 204140 101480 204360 101520
rect 204140 101410 204150 101480
rect 204350 101410 204360 101480
rect 204140 101360 204360 101410
rect 204640 101590 204860 101640
rect 204640 101520 204650 101590
rect 204850 101520 204860 101590
rect 204640 101480 204860 101520
rect 204640 101410 204650 101480
rect 204850 101410 204860 101480
rect 204640 101360 204860 101410
rect 205140 101590 205360 101640
rect 205140 101520 205150 101590
rect 205350 101520 205360 101590
rect 205140 101480 205360 101520
rect 205140 101410 205150 101480
rect 205350 101410 205360 101480
rect 205140 101360 205360 101410
rect 205640 101590 205860 101640
rect 205640 101520 205650 101590
rect 205850 101520 205860 101590
rect 205640 101480 205860 101520
rect 205640 101410 205650 101480
rect 205850 101410 205860 101480
rect 205640 101360 205860 101410
rect 206140 101590 206360 101640
rect 206140 101520 206150 101590
rect 206350 101520 206360 101590
rect 206140 101480 206360 101520
rect 206140 101410 206150 101480
rect 206350 101410 206360 101480
rect 206140 101360 206360 101410
rect 206640 101590 206860 101640
rect 206640 101520 206650 101590
rect 206850 101520 206860 101590
rect 206640 101480 206860 101520
rect 206640 101410 206650 101480
rect 206850 101410 206860 101480
rect 206640 101360 206860 101410
rect 207140 101590 207360 101640
rect 207140 101520 207150 101590
rect 207350 101520 207360 101590
rect 207140 101480 207360 101520
rect 207140 101410 207150 101480
rect 207350 101410 207360 101480
rect 207140 101360 207360 101410
rect 207640 101590 207860 101640
rect 207640 101520 207650 101590
rect 207850 101520 207860 101590
rect 207640 101480 207860 101520
rect 207640 101410 207650 101480
rect 207850 101410 207860 101480
rect 207640 101360 207860 101410
rect 196000 101350 208000 101360
rect 196000 101150 196020 101350
rect 196090 101150 196410 101350
rect 196480 101150 196520 101350
rect 196590 101150 196910 101350
rect 196980 101150 197020 101350
rect 197090 101150 197410 101350
rect 197480 101150 197520 101350
rect 197590 101150 197910 101350
rect 197980 101150 198020 101350
rect 198090 101150 198410 101350
rect 198480 101150 198520 101350
rect 198590 101150 198910 101350
rect 198980 101150 199020 101350
rect 199090 101150 199410 101350
rect 199480 101150 199520 101350
rect 199590 101150 199910 101350
rect 199980 101150 200020 101350
rect 200090 101150 200410 101350
rect 200480 101150 200520 101350
rect 200590 101150 200910 101350
rect 200980 101150 201020 101350
rect 201090 101150 201410 101350
rect 201480 101150 201520 101350
rect 201590 101150 201910 101350
rect 201980 101150 202020 101350
rect 202090 101150 202410 101350
rect 202480 101150 202520 101350
rect 202590 101150 202910 101350
rect 202980 101150 203020 101350
rect 203090 101150 203410 101350
rect 203480 101150 203520 101350
rect 203590 101150 203910 101350
rect 203980 101150 204020 101350
rect 204090 101150 204410 101350
rect 204480 101150 204520 101350
rect 204590 101150 204910 101350
rect 204980 101150 205020 101350
rect 205090 101150 205410 101350
rect 205480 101150 205520 101350
rect 205590 101150 205910 101350
rect 205980 101150 206020 101350
rect 206090 101150 206410 101350
rect 206480 101150 206520 101350
rect 206590 101150 206910 101350
rect 206980 101150 207020 101350
rect 207090 101150 207410 101350
rect 207480 101150 207520 101350
rect 207590 101150 207910 101350
rect 207980 101150 208000 101350
rect 196000 101140 208000 101150
rect 196140 101090 196360 101140
rect 196140 101020 196150 101090
rect 196350 101020 196360 101090
rect 196140 100980 196360 101020
rect 196140 100910 196150 100980
rect 196350 100910 196360 100980
rect 196140 100860 196360 100910
rect 196640 101090 196860 101140
rect 196640 101020 196650 101090
rect 196850 101020 196860 101090
rect 196640 100980 196860 101020
rect 196640 100910 196650 100980
rect 196850 100910 196860 100980
rect 196640 100860 196860 100910
rect 197140 101090 197360 101140
rect 197140 101020 197150 101090
rect 197350 101020 197360 101090
rect 197140 100980 197360 101020
rect 197140 100910 197150 100980
rect 197350 100910 197360 100980
rect 197140 100860 197360 100910
rect 197640 101090 197860 101140
rect 197640 101020 197650 101090
rect 197850 101020 197860 101090
rect 197640 100980 197860 101020
rect 197640 100910 197650 100980
rect 197850 100910 197860 100980
rect 197640 100860 197860 100910
rect 198140 101090 198360 101140
rect 198140 101020 198150 101090
rect 198350 101020 198360 101090
rect 198140 100980 198360 101020
rect 198140 100910 198150 100980
rect 198350 100910 198360 100980
rect 198140 100860 198360 100910
rect 198640 101090 198860 101140
rect 198640 101020 198650 101090
rect 198850 101020 198860 101090
rect 198640 100980 198860 101020
rect 198640 100910 198650 100980
rect 198850 100910 198860 100980
rect 198640 100860 198860 100910
rect 199140 101090 199360 101140
rect 199140 101020 199150 101090
rect 199350 101020 199360 101090
rect 199140 100980 199360 101020
rect 199140 100910 199150 100980
rect 199350 100910 199360 100980
rect 199140 100860 199360 100910
rect 199640 101090 199860 101140
rect 199640 101020 199650 101090
rect 199850 101020 199860 101090
rect 199640 100980 199860 101020
rect 199640 100910 199650 100980
rect 199850 100910 199860 100980
rect 199640 100860 199860 100910
rect 200140 101090 200360 101140
rect 200140 101020 200150 101090
rect 200350 101020 200360 101090
rect 200140 100980 200360 101020
rect 200140 100910 200150 100980
rect 200350 100910 200360 100980
rect 200140 100860 200360 100910
rect 200640 101090 200860 101140
rect 200640 101020 200650 101090
rect 200850 101020 200860 101090
rect 200640 100980 200860 101020
rect 200640 100910 200650 100980
rect 200850 100910 200860 100980
rect 200640 100860 200860 100910
rect 201140 101090 201360 101140
rect 201140 101020 201150 101090
rect 201350 101020 201360 101090
rect 201140 100980 201360 101020
rect 201140 100910 201150 100980
rect 201350 100910 201360 100980
rect 201140 100860 201360 100910
rect 201640 101090 201860 101140
rect 201640 101020 201650 101090
rect 201850 101020 201860 101090
rect 201640 100980 201860 101020
rect 201640 100910 201650 100980
rect 201850 100910 201860 100980
rect 201640 100860 201860 100910
rect 202140 101090 202360 101140
rect 202140 101020 202150 101090
rect 202350 101020 202360 101090
rect 202140 100980 202360 101020
rect 202140 100910 202150 100980
rect 202350 100910 202360 100980
rect 202140 100860 202360 100910
rect 202640 101090 202860 101140
rect 202640 101020 202650 101090
rect 202850 101020 202860 101090
rect 202640 100980 202860 101020
rect 202640 100910 202650 100980
rect 202850 100910 202860 100980
rect 202640 100860 202860 100910
rect 203140 101090 203360 101140
rect 203140 101020 203150 101090
rect 203350 101020 203360 101090
rect 203140 100980 203360 101020
rect 203140 100910 203150 100980
rect 203350 100910 203360 100980
rect 203140 100860 203360 100910
rect 203640 101090 203860 101140
rect 203640 101020 203650 101090
rect 203850 101020 203860 101090
rect 203640 100980 203860 101020
rect 203640 100910 203650 100980
rect 203850 100910 203860 100980
rect 203640 100860 203860 100910
rect 204140 101090 204360 101140
rect 204140 101020 204150 101090
rect 204350 101020 204360 101090
rect 204140 100980 204360 101020
rect 204140 100910 204150 100980
rect 204350 100910 204360 100980
rect 204140 100860 204360 100910
rect 204640 101090 204860 101140
rect 204640 101020 204650 101090
rect 204850 101020 204860 101090
rect 204640 100980 204860 101020
rect 204640 100910 204650 100980
rect 204850 100910 204860 100980
rect 204640 100860 204860 100910
rect 205140 101090 205360 101140
rect 205140 101020 205150 101090
rect 205350 101020 205360 101090
rect 205140 100980 205360 101020
rect 205140 100910 205150 100980
rect 205350 100910 205360 100980
rect 205140 100860 205360 100910
rect 205640 101090 205860 101140
rect 205640 101020 205650 101090
rect 205850 101020 205860 101090
rect 205640 100980 205860 101020
rect 205640 100910 205650 100980
rect 205850 100910 205860 100980
rect 205640 100860 205860 100910
rect 206140 101090 206360 101140
rect 206140 101020 206150 101090
rect 206350 101020 206360 101090
rect 206140 100980 206360 101020
rect 206140 100910 206150 100980
rect 206350 100910 206360 100980
rect 206140 100860 206360 100910
rect 206640 101090 206860 101140
rect 206640 101020 206650 101090
rect 206850 101020 206860 101090
rect 206640 100980 206860 101020
rect 206640 100910 206650 100980
rect 206850 100910 206860 100980
rect 206640 100860 206860 100910
rect 207140 101090 207360 101140
rect 207140 101020 207150 101090
rect 207350 101020 207360 101090
rect 207140 100980 207360 101020
rect 207140 100910 207150 100980
rect 207350 100910 207360 100980
rect 207140 100860 207360 100910
rect 207640 101090 207860 101140
rect 207640 101020 207650 101090
rect 207850 101020 207860 101090
rect 207640 100980 207860 101020
rect 207640 100910 207650 100980
rect 207850 100910 207860 100980
rect 207640 100860 207860 100910
rect 196000 100850 208000 100860
rect 196000 100650 196020 100850
rect 196090 100650 196410 100850
rect 196480 100650 196520 100850
rect 196590 100650 196910 100850
rect 196980 100650 197020 100850
rect 197090 100650 197410 100850
rect 197480 100650 197520 100850
rect 197590 100650 197910 100850
rect 197980 100650 198020 100850
rect 198090 100650 198410 100850
rect 198480 100650 198520 100850
rect 198590 100650 198910 100850
rect 198980 100650 199020 100850
rect 199090 100650 199410 100850
rect 199480 100650 199520 100850
rect 199590 100650 199910 100850
rect 199980 100650 200020 100850
rect 200090 100650 200410 100850
rect 200480 100650 200520 100850
rect 200590 100650 200910 100850
rect 200980 100650 201020 100850
rect 201090 100650 201410 100850
rect 201480 100650 201520 100850
rect 201590 100650 201910 100850
rect 201980 100650 202020 100850
rect 202090 100650 202410 100850
rect 202480 100650 202520 100850
rect 202590 100650 202910 100850
rect 202980 100650 203020 100850
rect 203090 100650 203410 100850
rect 203480 100650 203520 100850
rect 203590 100650 203910 100850
rect 203980 100650 204020 100850
rect 204090 100650 204410 100850
rect 204480 100650 204520 100850
rect 204590 100650 204910 100850
rect 204980 100650 205020 100850
rect 205090 100650 205410 100850
rect 205480 100650 205520 100850
rect 205590 100650 205910 100850
rect 205980 100650 206020 100850
rect 206090 100650 206410 100850
rect 206480 100650 206520 100850
rect 206590 100650 206910 100850
rect 206980 100650 207020 100850
rect 207090 100650 207410 100850
rect 207480 100650 207520 100850
rect 207590 100650 207910 100850
rect 207980 100650 208000 100850
rect 196000 100640 208000 100650
rect 196140 100590 196360 100640
rect 196140 100520 196150 100590
rect 196350 100520 196360 100590
rect 196140 100480 196360 100520
rect 196140 100410 196150 100480
rect 196350 100410 196360 100480
rect 196140 100360 196360 100410
rect 196640 100590 196860 100640
rect 196640 100520 196650 100590
rect 196850 100520 196860 100590
rect 196640 100480 196860 100520
rect 196640 100410 196650 100480
rect 196850 100410 196860 100480
rect 196640 100360 196860 100410
rect 197140 100590 197360 100640
rect 197140 100520 197150 100590
rect 197350 100520 197360 100590
rect 197140 100480 197360 100520
rect 197140 100410 197150 100480
rect 197350 100410 197360 100480
rect 197140 100360 197360 100410
rect 197640 100590 197860 100640
rect 197640 100520 197650 100590
rect 197850 100520 197860 100590
rect 197640 100480 197860 100520
rect 197640 100410 197650 100480
rect 197850 100410 197860 100480
rect 197640 100360 197860 100410
rect 198140 100590 198360 100640
rect 198140 100520 198150 100590
rect 198350 100520 198360 100590
rect 198140 100480 198360 100520
rect 198140 100410 198150 100480
rect 198350 100410 198360 100480
rect 198140 100360 198360 100410
rect 198640 100590 198860 100640
rect 198640 100520 198650 100590
rect 198850 100520 198860 100590
rect 198640 100480 198860 100520
rect 198640 100410 198650 100480
rect 198850 100410 198860 100480
rect 198640 100360 198860 100410
rect 199140 100590 199360 100640
rect 199140 100520 199150 100590
rect 199350 100520 199360 100590
rect 199140 100480 199360 100520
rect 199140 100410 199150 100480
rect 199350 100410 199360 100480
rect 199140 100360 199360 100410
rect 199640 100590 199860 100640
rect 199640 100520 199650 100590
rect 199850 100520 199860 100590
rect 199640 100480 199860 100520
rect 199640 100410 199650 100480
rect 199850 100410 199860 100480
rect 199640 100360 199860 100410
rect 200140 100590 200360 100640
rect 200140 100520 200150 100590
rect 200350 100520 200360 100590
rect 200140 100480 200360 100520
rect 200140 100410 200150 100480
rect 200350 100410 200360 100480
rect 200140 100360 200360 100410
rect 200640 100590 200860 100640
rect 200640 100520 200650 100590
rect 200850 100520 200860 100590
rect 200640 100480 200860 100520
rect 200640 100410 200650 100480
rect 200850 100410 200860 100480
rect 200640 100360 200860 100410
rect 201140 100590 201360 100640
rect 201140 100520 201150 100590
rect 201350 100520 201360 100590
rect 201140 100480 201360 100520
rect 201140 100410 201150 100480
rect 201350 100410 201360 100480
rect 201140 100360 201360 100410
rect 201640 100590 201860 100640
rect 201640 100520 201650 100590
rect 201850 100520 201860 100590
rect 201640 100480 201860 100520
rect 201640 100410 201650 100480
rect 201850 100410 201860 100480
rect 201640 100360 201860 100410
rect 202140 100590 202360 100640
rect 202140 100520 202150 100590
rect 202350 100520 202360 100590
rect 202140 100480 202360 100520
rect 202140 100410 202150 100480
rect 202350 100410 202360 100480
rect 202140 100360 202360 100410
rect 202640 100590 202860 100640
rect 202640 100520 202650 100590
rect 202850 100520 202860 100590
rect 202640 100480 202860 100520
rect 202640 100410 202650 100480
rect 202850 100410 202860 100480
rect 202640 100360 202860 100410
rect 203140 100590 203360 100640
rect 203140 100520 203150 100590
rect 203350 100520 203360 100590
rect 203140 100480 203360 100520
rect 203140 100410 203150 100480
rect 203350 100410 203360 100480
rect 203140 100360 203360 100410
rect 203640 100590 203860 100640
rect 203640 100520 203650 100590
rect 203850 100520 203860 100590
rect 203640 100480 203860 100520
rect 203640 100410 203650 100480
rect 203850 100410 203860 100480
rect 203640 100360 203860 100410
rect 204140 100590 204360 100640
rect 204140 100520 204150 100590
rect 204350 100520 204360 100590
rect 204140 100480 204360 100520
rect 204140 100410 204150 100480
rect 204350 100410 204360 100480
rect 204140 100360 204360 100410
rect 204640 100590 204860 100640
rect 204640 100520 204650 100590
rect 204850 100520 204860 100590
rect 204640 100480 204860 100520
rect 204640 100410 204650 100480
rect 204850 100410 204860 100480
rect 204640 100360 204860 100410
rect 205140 100590 205360 100640
rect 205140 100520 205150 100590
rect 205350 100520 205360 100590
rect 205140 100480 205360 100520
rect 205140 100410 205150 100480
rect 205350 100410 205360 100480
rect 205140 100360 205360 100410
rect 205640 100590 205860 100640
rect 205640 100520 205650 100590
rect 205850 100520 205860 100590
rect 205640 100480 205860 100520
rect 205640 100410 205650 100480
rect 205850 100410 205860 100480
rect 205640 100360 205860 100410
rect 206140 100590 206360 100640
rect 206140 100520 206150 100590
rect 206350 100520 206360 100590
rect 206140 100480 206360 100520
rect 206140 100410 206150 100480
rect 206350 100410 206360 100480
rect 206140 100360 206360 100410
rect 206640 100590 206860 100640
rect 206640 100520 206650 100590
rect 206850 100520 206860 100590
rect 206640 100480 206860 100520
rect 206640 100410 206650 100480
rect 206850 100410 206860 100480
rect 206640 100360 206860 100410
rect 207140 100590 207360 100640
rect 207140 100520 207150 100590
rect 207350 100520 207360 100590
rect 207140 100480 207360 100520
rect 207140 100410 207150 100480
rect 207350 100410 207360 100480
rect 207140 100360 207360 100410
rect 207640 100590 207860 100640
rect 207640 100520 207650 100590
rect 207850 100520 207860 100590
rect 207640 100480 207860 100520
rect 207640 100410 207650 100480
rect 207850 100410 207860 100480
rect 207640 100360 207860 100410
rect 196000 100350 208000 100360
rect 196000 100150 196020 100350
rect 196090 100150 196410 100350
rect 196480 100150 196520 100350
rect 196590 100150 196910 100350
rect 196980 100150 197020 100350
rect 197090 100150 197410 100350
rect 197480 100150 197520 100350
rect 197590 100150 197910 100350
rect 197980 100150 198020 100350
rect 198090 100150 198410 100350
rect 198480 100150 198520 100350
rect 198590 100150 198910 100350
rect 198980 100150 199020 100350
rect 199090 100150 199410 100350
rect 199480 100150 199520 100350
rect 199590 100150 199910 100350
rect 199980 100150 200020 100350
rect 200090 100150 200410 100350
rect 200480 100150 200520 100350
rect 200590 100150 200910 100350
rect 200980 100150 201020 100350
rect 201090 100150 201410 100350
rect 201480 100150 201520 100350
rect 201590 100150 201910 100350
rect 201980 100150 202020 100350
rect 202090 100150 202410 100350
rect 202480 100150 202520 100350
rect 202590 100150 202910 100350
rect 202980 100150 203020 100350
rect 203090 100150 203410 100350
rect 203480 100150 203520 100350
rect 203590 100150 203910 100350
rect 203980 100150 204020 100350
rect 204090 100150 204410 100350
rect 204480 100150 204520 100350
rect 204590 100150 204910 100350
rect 204980 100150 205020 100350
rect 205090 100150 205410 100350
rect 205480 100150 205520 100350
rect 205590 100150 205910 100350
rect 205980 100150 206020 100350
rect 206090 100150 206410 100350
rect 206480 100150 206520 100350
rect 206590 100150 206910 100350
rect 206980 100150 207020 100350
rect 207090 100150 207410 100350
rect 207480 100150 207520 100350
rect 207590 100150 207910 100350
rect 207980 100150 208000 100350
rect 196000 100140 208000 100150
rect 196140 100090 196360 100140
rect 196140 100020 196150 100090
rect 196350 100020 196360 100090
rect 196140 99980 196360 100020
rect 196140 99910 196150 99980
rect 196350 99910 196360 99980
rect 196140 99860 196360 99910
rect 196640 100090 196860 100140
rect 196640 100020 196650 100090
rect 196850 100020 196860 100090
rect 196640 99980 196860 100020
rect 196640 99910 196650 99980
rect 196850 99910 196860 99980
rect 196640 99860 196860 99910
rect 197140 100090 197360 100140
rect 197140 100020 197150 100090
rect 197350 100020 197360 100090
rect 197140 99980 197360 100020
rect 197140 99910 197150 99980
rect 197350 99910 197360 99980
rect 197140 99860 197360 99910
rect 197640 100090 197860 100140
rect 197640 100020 197650 100090
rect 197850 100020 197860 100090
rect 197640 99980 197860 100020
rect 197640 99910 197650 99980
rect 197850 99910 197860 99980
rect 197640 99860 197860 99910
rect 198140 100090 198360 100140
rect 198140 100020 198150 100090
rect 198350 100020 198360 100090
rect 198140 99980 198360 100020
rect 198140 99910 198150 99980
rect 198350 99910 198360 99980
rect 198140 99860 198360 99910
rect 198640 100090 198860 100140
rect 198640 100020 198650 100090
rect 198850 100020 198860 100090
rect 198640 99980 198860 100020
rect 198640 99910 198650 99980
rect 198850 99910 198860 99980
rect 198640 99860 198860 99910
rect 199140 100090 199360 100140
rect 199140 100020 199150 100090
rect 199350 100020 199360 100090
rect 199140 99980 199360 100020
rect 199140 99910 199150 99980
rect 199350 99910 199360 99980
rect 199140 99860 199360 99910
rect 199640 100090 199860 100140
rect 199640 100020 199650 100090
rect 199850 100020 199860 100090
rect 199640 99980 199860 100020
rect 199640 99910 199650 99980
rect 199850 99910 199860 99980
rect 199640 99860 199860 99910
rect 200140 100090 200360 100140
rect 200140 100020 200150 100090
rect 200350 100020 200360 100090
rect 200140 99980 200360 100020
rect 200140 99910 200150 99980
rect 200350 99910 200360 99980
rect 200140 99860 200360 99910
rect 200640 100090 200860 100140
rect 200640 100020 200650 100090
rect 200850 100020 200860 100090
rect 200640 99980 200860 100020
rect 200640 99910 200650 99980
rect 200850 99910 200860 99980
rect 200640 99860 200860 99910
rect 201140 100090 201360 100140
rect 201140 100020 201150 100090
rect 201350 100020 201360 100090
rect 201140 99980 201360 100020
rect 201140 99910 201150 99980
rect 201350 99910 201360 99980
rect 201140 99860 201360 99910
rect 201640 100090 201860 100140
rect 201640 100020 201650 100090
rect 201850 100020 201860 100090
rect 201640 99980 201860 100020
rect 201640 99910 201650 99980
rect 201850 99910 201860 99980
rect 201640 99860 201860 99910
rect 202140 100090 202360 100140
rect 202140 100020 202150 100090
rect 202350 100020 202360 100090
rect 202140 99980 202360 100020
rect 202140 99910 202150 99980
rect 202350 99910 202360 99980
rect 202140 99860 202360 99910
rect 202640 100090 202860 100140
rect 202640 100020 202650 100090
rect 202850 100020 202860 100090
rect 202640 99980 202860 100020
rect 202640 99910 202650 99980
rect 202850 99910 202860 99980
rect 202640 99860 202860 99910
rect 203140 100090 203360 100140
rect 203140 100020 203150 100090
rect 203350 100020 203360 100090
rect 203140 99980 203360 100020
rect 203140 99910 203150 99980
rect 203350 99910 203360 99980
rect 203140 99860 203360 99910
rect 203640 100090 203860 100140
rect 203640 100020 203650 100090
rect 203850 100020 203860 100090
rect 203640 99980 203860 100020
rect 203640 99910 203650 99980
rect 203850 99910 203860 99980
rect 203640 99860 203860 99910
rect 204140 100090 204360 100140
rect 204140 100020 204150 100090
rect 204350 100020 204360 100090
rect 204140 99980 204360 100020
rect 204140 99910 204150 99980
rect 204350 99910 204360 99980
rect 204140 99860 204360 99910
rect 204640 100090 204860 100140
rect 204640 100020 204650 100090
rect 204850 100020 204860 100090
rect 204640 99980 204860 100020
rect 204640 99910 204650 99980
rect 204850 99910 204860 99980
rect 204640 99860 204860 99910
rect 205140 100090 205360 100140
rect 205140 100020 205150 100090
rect 205350 100020 205360 100090
rect 205140 99980 205360 100020
rect 205140 99910 205150 99980
rect 205350 99910 205360 99980
rect 205140 99860 205360 99910
rect 205640 100090 205860 100140
rect 205640 100020 205650 100090
rect 205850 100020 205860 100090
rect 205640 99980 205860 100020
rect 205640 99910 205650 99980
rect 205850 99910 205860 99980
rect 205640 99860 205860 99910
rect 206140 100090 206360 100140
rect 206140 100020 206150 100090
rect 206350 100020 206360 100090
rect 206140 99980 206360 100020
rect 206140 99910 206150 99980
rect 206350 99910 206360 99980
rect 206140 99860 206360 99910
rect 206640 100090 206860 100140
rect 206640 100020 206650 100090
rect 206850 100020 206860 100090
rect 206640 99980 206860 100020
rect 206640 99910 206650 99980
rect 206850 99910 206860 99980
rect 206640 99860 206860 99910
rect 207140 100090 207360 100140
rect 207140 100020 207150 100090
rect 207350 100020 207360 100090
rect 207140 99980 207360 100020
rect 207140 99910 207150 99980
rect 207350 99910 207360 99980
rect 207140 99860 207360 99910
rect 207640 100090 207860 100140
rect 207640 100020 207650 100090
rect 207850 100020 207860 100090
rect 207640 99980 207860 100020
rect 207640 99910 207650 99980
rect 207850 99910 207860 99980
rect 207640 99860 207860 99910
rect 196000 99850 208000 99860
rect 196000 99650 196020 99850
rect 196090 99650 196410 99850
rect 196480 99650 196520 99850
rect 196590 99650 196910 99850
rect 196980 99650 197020 99850
rect 197090 99650 197410 99850
rect 197480 99650 197520 99850
rect 197590 99650 197910 99850
rect 197980 99650 198020 99850
rect 198090 99650 198410 99850
rect 198480 99650 198520 99850
rect 198590 99650 198910 99850
rect 198980 99650 199020 99850
rect 199090 99650 199410 99850
rect 199480 99650 199520 99850
rect 199590 99650 199910 99850
rect 199980 99650 200020 99850
rect 200090 99650 200410 99850
rect 200480 99650 200520 99850
rect 200590 99650 200910 99850
rect 200980 99650 201020 99850
rect 201090 99650 201410 99850
rect 201480 99650 201520 99850
rect 201590 99650 201910 99850
rect 201980 99650 202020 99850
rect 202090 99650 202410 99850
rect 202480 99650 202520 99850
rect 202590 99650 202910 99850
rect 202980 99650 203020 99850
rect 203090 99650 203410 99850
rect 203480 99650 203520 99850
rect 203590 99650 203910 99850
rect 203980 99650 204020 99850
rect 204090 99650 204410 99850
rect 204480 99650 204520 99850
rect 204590 99650 204910 99850
rect 204980 99650 205020 99850
rect 205090 99650 205410 99850
rect 205480 99650 205520 99850
rect 205590 99650 205910 99850
rect 205980 99650 206020 99850
rect 206090 99650 206410 99850
rect 206480 99650 206520 99850
rect 206590 99650 206910 99850
rect 206980 99650 207020 99850
rect 207090 99650 207410 99850
rect 207480 99650 207520 99850
rect 207590 99650 207910 99850
rect 207980 99650 208000 99850
rect 196000 99640 208000 99650
rect 196140 99590 196360 99640
rect 196140 99520 196150 99590
rect 196350 99520 196360 99590
rect 196140 99480 196360 99520
rect 196140 99410 196150 99480
rect 196350 99410 196360 99480
rect 196140 99360 196360 99410
rect 196640 99590 196860 99640
rect 196640 99520 196650 99590
rect 196850 99520 196860 99590
rect 196640 99480 196860 99520
rect 196640 99410 196650 99480
rect 196850 99410 196860 99480
rect 196640 99360 196860 99410
rect 197140 99590 197360 99640
rect 197140 99520 197150 99590
rect 197350 99520 197360 99590
rect 197140 99480 197360 99520
rect 197140 99410 197150 99480
rect 197350 99410 197360 99480
rect 197140 99360 197360 99410
rect 197640 99590 197860 99640
rect 197640 99520 197650 99590
rect 197850 99520 197860 99590
rect 197640 99480 197860 99520
rect 197640 99410 197650 99480
rect 197850 99410 197860 99480
rect 197640 99360 197860 99410
rect 198140 99590 198360 99640
rect 198140 99520 198150 99590
rect 198350 99520 198360 99590
rect 198140 99480 198360 99520
rect 198140 99410 198150 99480
rect 198350 99410 198360 99480
rect 198140 99360 198360 99410
rect 198640 99590 198860 99640
rect 198640 99520 198650 99590
rect 198850 99520 198860 99590
rect 198640 99480 198860 99520
rect 198640 99410 198650 99480
rect 198850 99410 198860 99480
rect 198640 99360 198860 99410
rect 199140 99590 199360 99640
rect 199140 99520 199150 99590
rect 199350 99520 199360 99590
rect 199140 99480 199360 99520
rect 199140 99410 199150 99480
rect 199350 99410 199360 99480
rect 199140 99360 199360 99410
rect 199640 99590 199860 99640
rect 199640 99520 199650 99590
rect 199850 99520 199860 99590
rect 199640 99480 199860 99520
rect 199640 99410 199650 99480
rect 199850 99410 199860 99480
rect 199640 99360 199860 99410
rect 200140 99590 200360 99640
rect 200140 99520 200150 99590
rect 200350 99520 200360 99590
rect 200140 99480 200360 99520
rect 200140 99410 200150 99480
rect 200350 99410 200360 99480
rect 200140 99360 200360 99410
rect 200640 99590 200860 99640
rect 200640 99520 200650 99590
rect 200850 99520 200860 99590
rect 200640 99480 200860 99520
rect 200640 99410 200650 99480
rect 200850 99410 200860 99480
rect 200640 99360 200860 99410
rect 201140 99590 201360 99640
rect 201140 99520 201150 99590
rect 201350 99520 201360 99590
rect 201140 99480 201360 99520
rect 201140 99410 201150 99480
rect 201350 99410 201360 99480
rect 201140 99360 201360 99410
rect 201640 99590 201860 99640
rect 201640 99520 201650 99590
rect 201850 99520 201860 99590
rect 201640 99480 201860 99520
rect 201640 99410 201650 99480
rect 201850 99410 201860 99480
rect 201640 99360 201860 99410
rect 202140 99590 202360 99640
rect 202140 99520 202150 99590
rect 202350 99520 202360 99590
rect 202140 99480 202360 99520
rect 202140 99410 202150 99480
rect 202350 99410 202360 99480
rect 202140 99360 202360 99410
rect 202640 99590 202860 99640
rect 202640 99520 202650 99590
rect 202850 99520 202860 99590
rect 202640 99480 202860 99520
rect 202640 99410 202650 99480
rect 202850 99410 202860 99480
rect 202640 99360 202860 99410
rect 203140 99590 203360 99640
rect 203140 99520 203150 99590
rect 203350 99520 203360 99590
rect 203140 99480 203360 99520
rect 203140 99410 203150 99480
rect 203350 99410 203360 99480
rect 203140 99360 203360 99410
rect 203640 99590 203860 99640
rect 203640 99520 203650 99590
rect 203850 99520 203860 99590
rect 203640 99480 203860 99520
rect 203640 99410 203650 99480
rect 203850 99410 203860 99480
rect 203640 99360 203860 99410
rect 204140 99590 204360 99640
rect 204140 99520 204150 99590
rect 204350 99520 204360 99590
rect 204140 99480 204360 99520
rect 204140 99410 204150 99480
rect 204350 99410 204360 99480
rect 204140 99360 204360 99410
rect 204640 99590 204860 99640
rect 204640 99520 204650 99590
rect 204850 99520 204860 99590
rect 204640 99480 204860 99520
rect 204640 99410 204650 99480
rect 204850 99410 204860 99480
rect 204640 99360 204860 99410
rect 205140 99590 205360 99640
rect 205140 99520 205150 99590
rect 205350 99520 205360 99590
rect 205140 99480 205360 99520
rect 205140 99410 205150 99480
rect 205350 99410 205360 99480
rect 205140 99360 205360 99410
rect 205640 99590 205860 99640
rect 205640 99520 205650 99590
rect 205850 99520 205860 99590
rect 205640 99480 205860 99520
rect 205640 99410 205650 99480
rect 205850 99410 205860 99480
rect 205640 99360 205860 99410
rect 206140 99590 206360 99640
rect 206140 99520 206150 99590
rect 206350 99520 206360 99590
rect 206140 99480 206360 99520
rect 206140 99410 206150 99480
rect 206350 99410 206360 99480
rect 206140 99360 206360 99410
rect 206640 99590 206860 99640
rect 206640 99520 206650 99590
rect 206850 99520 206860 99590
rect 206640 99480 206860 99520
rect 206640 99410 206650 99480
rect 206850 99410 206860 99480
rect 206640 99360 206860 99410
rect 207140 99590 207360 99640
rect 207140 99520 207150 99590
rect 207350 99520 207360 99590
rect 207140 99480 207360 99520
rect 207140 99410 207150 99480
rect 207350 99410 207360 99480
rect 207140 99360 207360 99410
rect 207640 99590 207860 99640
rect 207640 99520 207650 99590
rect 207850 99520 207860 99590
rect 207640 99480 207860 99520
rect 207640 99410 207650 99480
rect 207850 99410 207860 99480
rect 207640 99360 207860 99410
rect 196000 99350 208000 99360
rect 196000 99150 196020 99350
rect 196090 99150 196410 99350
rect 196480 99150 196520 99350
rect 196590 99150 196910 99350
rect 196980 99150 197020 99350
rect 197090 99150 197410 99350
rect 197480 99150 197520 99350
rect 197590 99150 197910 99350
rect 197980 99150 198020 99350
rect 198090 99150 198410 99350
rect 198480 99150 198520 99350
rect 198590 99150 198910 99350
rect 198980 99150 199020 99350
rect 199090 99150 199410 99350
rect 199480 99150 199520 99350
rect 199590 99150 199910 99350
rect 199980 99150 200020 99350
rect 200090 99150 200410 99350
rect 200480 99150 200520 99350
rect 200590 99150 200910 99350
rect 200980 99150 201020 99350
rect 201090 99150 201410 99350
rect 201480 99150 201520 99350
rect 201590 99150 201910 99350
rect 201980 99150 202020 99350
rect 202090 99150 202410 99350
rect 202480 99150 202520 99350
rect 202590 99150 202910 99350
rect 202980 99150 203020 99350
rect 203090 99150 203410 99350
rect 203480 99150 203520 99350
rect 203590 99150 203910 99350
rect 203980 99150 204020 99350
rect 204090 99150 204410 99350
rect 204480 99150 204520 99350
rect 204590 99150 204910 99350
rect 204980 99150 205020 99350
rect 205090 99150 205410 99350
rect 205480 99150 205520 99350
rect 205590 99150 205910 99350
rect 205980 99150 206020 99350
rect 206090 99150 206410 99350
rect 206480 99150 206520 99350
rect 206590 99150 206910 99350
rect 206980 99150 207020 99350
rect 207090 99150 207410 99350
rect 207480 99150 207520 99350
rect 207590 99150 207910 99350
rect 207980 99150 208000 99350
rect 196000 99140 208000 99150
rect 196140 99090 196360 99140
rect 196140 99020 196150 99090
rect 196350 99020 196360 99090
rect 196140 98980 196360 99020
rect 196140 98910 196150 98980
rect 196350 98910 196360 98980
rect 196140 98860 196360 98910
rect 196640 99090 196860 99140
rect 196640 99020 196650 99090
rect 196850 99020 196860 99090
rect 196640 98980 196860 99020
rect 196640 98910 196650 98980
rect 196850 98910 196860 98980
rect 196640 98860 196860 98910
rect 197140 99090 197360 99140
rect 197140 99020 197150 99090
rect 197350 99020 197360 99090
rect 197140 98980 197360 99020
rect 197140 98910 197150 98980
rect 197350 98910 197360 98980
rect 197140 98860 197360 98910
rect 197640 99090 197860 99140
rect 197640 99020 197650 99090
rect 197850 99020 197860 99090
rect 197640 98980 197860 99020
rect 197640 98910 197650 98980
rect 197850 98910 197860 98980
rect 197640 98860 197860 98910
rect 198140 99090 198360 99140
rect 198140 99020 198150 99090
rect 198350 99020 198360 99090
rect 198140 98980 198360 99020
rect 198140 98910 198150 98980
rect 198350 98910 198360 98980
rect 198140 98860 198360 98910
rect 198640 99090 198860 99140
rect 198640 99020 198650 99090
rect 198850 99020 198860 99090
rect 198640 98980 198860 99020
rect 198640 98910 198650 98980
rect 198850 98910 198860 98980
rect 198640 98860 198860 98910
rect 199140 99090 199360 99140
rect 199140 99020 199150 99090
rect 199350 99020 199360 99090
rect 199140 98980 199360 99020
rect 199140 98910 199150 98980
rect 199350 98910 199360 98980
rect 199140 98860 199360 98910
rect 199640 99090 199860 99140
rect 199640 99020 199650 99090
rect 199850 99020 199860 99090
rect 199640 98980 199860 99020
rect 199640 98910 199650 98980
rect 199850 98910 199860 98980
rect 199640 98860 199860 98910
rect 200140 99090 200360 99140
rect 200140 99020 200150 99090
rect 200350 99020 200360 99090
rect 200140 98980 200360 99020
rect 200140 98910 200150 98980
rect 200350 98910 200360 98980
rect 200140 98860 200360 98910
rect 200640 99090 200860 99140
rect 200640 99020 200650 99090
rect 200850 99020 200860 99090
rect 200640 98980 200860 99020
rect 200640 98910 200650 98980
rect 200850 98910 200860 98980
rect 200640 98860 200860 98910
rect 201140 99090 201360 99140
rect 201140 99020 201150 99090
rect 201350 99020 201360 99090
rect 201140 98980 201360 99020
rect 201140 98910 201150 98980
rect 201350 98910 201360 98980
rect 201140 98860 201360 98910
rect 201640 99090 201860 99140
rect 201640 99020 201650 99090
rect 201850 99020 201860 99090
rect 201640 98980 201860 99020
rect 201640 98910 201650 98980
rect 201850 98910 201860 98980
rect 201640 98860 201860 98910
rect 202140 99090 202360 99140
rect 202140 99020 202150 99090
rect 202350 99020 202360 99090
rect 202140 98980 202360 99020
rect 202140 98910 202150 98980
rect 202350 98910 202360 98980
rect 202140 98860 202360 98910
rect 202640 99090 202860 99140
rect 202640 99020 202650 99090
rect 202850 99020 202860 99090
rect 202640 98980 202860 99020
rect 202640 98910 202650 98980
rect 202850 98910 202860 98980
rect 202640 98860 202860 98910
rect 203140 99090 203360 99140
rect 203140 99020 203150 99090
rect 203350 99020 203360 99090
rect 203140 98980 203360 99020
rect 203140 98910 203150 98980
rect 203350 98910 203360 98980
rect 203140 98860 203360 98910
rect 203640 99090 203860 99140
rect 203640 99020 203650 99090
rect 203850 99020 203860 99090
rect 203640 98980 203860 99020
rect 203640 98910 203650 98980
rect 203850 98910 203860 98980
rect 203640 98860 203860 98910
rect 204140 99090 204360 99140
rect 204140 99020 204150 99090
rect 204350 99020 204360 99090
rect 204140 98980 204360 99020
rect 204140 98910 204150 98980
rect 204350 98910 204360 98980
rect 204140 98860 204360 98910
rect 204640 99090 204860 99140
rect 204640 99020 204650 99090
rect 204850 99020 204860 99090
rect 204640 98980 204860 99020
rect 204640 98910 204650 98980
rect 204850 98910 204860 98980
rect 204640 98860 204860 98910
rect 205140 99090 205360 99140
rect 205140 99020 205150 99090
rect 205350 99020 205360 99090
rect 205140 98980 205360 99020
rect 205140 98910 205150 98980
rect 205350 98910 205360 98980
rect 205140 98860 205360 98910
rect 205640 99090 205860 99140
rect 205640 99020 205650 99090
rect 205850 99020 205860 99090
rect 205640 98980 205860 99020
rect 205640 98910 205650 98980
rect 205850 98910 205860 98980
rect 205640 98860 205860 98910
rect 206140 99090 206360 99140
rect 206140 99020 206150 99090
rect 206350 99020 206360 99090
rect 206140 98980 206360 99020
rect 206140 98910 206150 98980
rect 206350 98910 206360 98980
rect 206140 98860 206360 98910
rect 206640 99090 206860 99140
rect 206640 99020 206650 99090
rect 206850 99020 206860 99090
rect 206640 98980 206860 99020
rect 206640 98910 206650 98980
rect 206850 98910 206860 98980
rect 206640 98860 206860 98910
rect 207140 99090 207360 99140
rect 207140 99020 207150 99090
rect 207350 99020 207360 99090
rect 207140 98980 207360 99020
rect 207140 98910 207150 98980
rect 207350 98910 207360 98980
rect 207140 98860 207360 98910
rect 207640 99090 207860 99140
rect 207640 99020 207650 99090
rect 207850 99020 207860 99090
rect 207640 98980 207860 99020
rect 207640 98910 207650 98980
rect 207850 98910 207860 98980
rect 207640 98860 207860 98910
rect 196000 98850 208000 98860
rect 196000 98650 196020 98850
rect 196090 98650 196410 98850
rect 196480 98650 196520 98850
rect 196590 98650 196910 98850
rect 196980 98650 197020 98850
rect 197090 98650 197410 98850
rect 197480 98650 197520 98850
rect 197590 98650 197910 98850
rect 197980 98650 198020 98850
rect 198090 98650 198410 98850
rect 198480 98650 198520 98850
rect 198590 98650 198910 98850
rect 198980 98650 199020 98850
rect 199090 98650 199410 98850
rect 199480 98650 199520 98850
rect 199590 98650 199910 98850
rect 199980 98650 200020 98850
rect 200090 98650 200410 98850
rect 200480 98650 200520 98850
rect 200590 98650 200910 98850
rect 200980 98650 201020 98850
rect 201090 98650 201410 98850
rect 201480 98650 201520 98850
rect 201590 98650 201910 98850
rect 201980 98650 202020 98850
rect 202090 98650 202410 98850
rect 202480 98650 202520 98850
rect 202590 98650 202910 98850
rect 202980 98650 203020 98850
rect 203090 98650 203410 98850
rect 203480 98650 203520 98850
rect 203590 98650 203910 98850
rect 203980 98650 204020 98850
rect 204090 98650 204410 98850
rect 204480 98650 204520 98850
rect 204590 98650 204910 98850
rect 204980 98650 205020 98850
rect 205090 98650 205410 98850
rect 205480 98650 205520 98850
rect 205590 98650 205910 98850
rect 205980 98650 206020 98850
rect 206090 98650 206410 98850
rect 206480 98650 206520 98850
rect 206590 98650 206910 98850
rect 206980 98650 207020 98850
rect 207090 98650 207410 98850
rect 207480 98650 207520 98850
rect 207590 98650 207910 98850
rect 207980 98650 208000 98850
rect 196000 98640 208000 98650
rect 196140 98590 196360 98640
rect 196140 98520 196150 98590
rect 196350 98520 196360 98590
rect 196140 98480 196360 98520
rect 196140 98410 196150 98480
rect 196350 98410 196360 98480
rect 196140 98360 196360 98410
rect 196640 98590 196860 98640
rect 196640 98520 196650 98590
rect 196850 98520 196860 98590
rect 196640 98480 196860 98520
rect 196640 98410 196650 98480
rect 196850 98410 196860 98480
rect 196640 98360 196860 98410
rect 197140 98590 197360 98640
rect 197140 98520 197150 98590
rect 197350 98520 197360 98590
rect 197140 98480 197360 98520
rect 197140 98410 197150 98480
rect 197350 98410 197360 98480
rect 197140 98360 197360 98410
rect 197640 98590 197860 98640
rect 197640 98520 197650 98590
rect 197850 98520 197860 98590
rect 197640 98480 197860 98520
rect 197640 98410 197650 98480
rect 197850 98410 197860 98480
rect 197640 98360 197860 98410
rect 198140 98590 198360 98640
rect 198140 98520 198150 98590
rect 198350 98520 198360 98590
rect 198140 98480 198360 98520
rect 198140 98410 198150 98480
rect 198350 98410 198360 98480
rect 198140 98360 198360 98410
rect 198640 98590 198860 98640
rect 198640 98520 198650 98590
rect 198850 98520 198860 98590
rect 198640 98480 198860 98520
rect 198640 98410 198650 98480
rect 198850 98410 198860 98480
rect 198640 98360 198860 98410
rect 199140 98590 199360 98640
rect 199140 98520 199150 98590
rect 199350 98520 199360 98590
rect 199140 98480 199360 98520
rect 199140 98410 199150 98480
rect 199350 98410 199360 98480
rect 199140 98360 199360 98410
rect 199640 98590 199860 98640
rect 199640 98520 199650 98590
rect 199850 98520 199860 98590
rect 199640 98480 199860 98520
rect 199640 98410 199650 98480
rect 199850 98410 199860 98480
rect 199640 98360 199860 98410
rect 200140 98590 200360 98640
rect 200140 98520 200150 98590
rect 200350 98520 200360 98590
rect 200140 98480 200360 98520
rect 200140 98410 200150 98480
rect 200350 98410 200360 98480
rect 200140 98360 200360 98410
rect 200640 98590 200860 98640
rect 200640 98520 200650 98590
rect 200850 98520 200860 98590
rect 200640 98480 200860 98520
rect 200640 98410 200650 98480
rect 200850 98410 200860 98480
rect 200640 98360 200860 98410
rect 201140 98590 201360 98640
rect 201140 98520 201150 98590
rect 201350 98520 201360 98590
rect 201140 98480 201360 98520
rect 201140 98410 201150 98480
rect 201350 98410 201360 98480
rect 201140 98360 201360 98410
rect 201640 98590 201860 98640
rect 201640 98520 201650 98590
rect 201850 98520 201860 98590
rect 201640 98480 201860 98520
rect 201640 98410 201650 98480
rect 201850 98410 201860 98480
rect 201640 98360 201860 98410
rect 202140 98590 202360 98640
rect 202140 98520 202150 98590
rect 202350 98520 202360 98590
rect 202140 98480 202360 98520
rect 202140 98410 202150 98480
rect 202350 98410 202360 98480
rect 202140 98360 202360 98410
rect 202640 98590 202860 98640
rect 202640 98520 202650 98590
rect 202850 98520 202860 98590
rect 202640 98480 202860 98520
rect 202640 98410 202650 98480
rect 202850 98410 202860 98480
rect 202640 98360 202860 98410
rect 203140 98590 203360 98640
rect 203140 98520 203150 98590
rect 203350 98520 203360 98590
rect 203140 98480 203360 98520
rect 203140 98410 203150 98480
rect 203350 98410 203360 98480
rect 203140 98360 203360 98410
rect 203640 98590 203860 98640
rect 203640 98520 203650 98590
rect 203850 98520 203860 98590
rect 203640 98480 203860 98520
rect 203640 98410 203650 98480
rect 203850 98410 203860 98480
rect 203640 98360 203860 98410
rect 204140 98590 204360 98640
rect 204140 98520 204150 98590
rect 204350 98520 204360 98590
rect 204140 98480 204360 98520
rect 204140 98410 204150 98480
rect 204350 98410 204360 98480
rect 204140 98360 204360 98410
rect 204640 98590 204860 98640
rect 204640 98520 204650 98590
rect 204850 98520 204860 98590
rect 204640 98480 204860 98520
rect 204640 98410 204650 98480
rect 204850 98410 204860 98480
rect 204640 98360 204860 98410
rect 205140 98590 205360 98640
rect 205140 98520 205150 98590
rect 205350 98520 205360 98590
rect 205140 98480 205360 98520
rect 205140 98410 205150 98480
rect 205350 98410 205360 98480
rect 205140 98360 205360 98410
rect 205640 98590 205860 98640
rect 205640 98520 205650 98590
rect 205850 98520 205860 98590
rect 205640 98480 205860 98520
rect 205640 98410 205650 98480
rect 205850 98410 205860 98480
rect 205640 98360 205860 98410
rect 206140 98590 206360 98640
rect 206140 98520 206150 98590
rect 206350 98520 206360 98590
rect 206140 98480 206360 98520
rect 206140 98410 206150 98480
rect 206350 98410 206360 98480
rect 206140 98360 206360 98410
rect 206640 98590 206860 98640
rect 206640 98520 206650 98590
rect 206850 98520 206860 98590
rect 206640 98480 206860 98520
rect 206640 98410 206650 98480
rect 206850 98410 206860 98480
rect 206640 98360 206860 98410
rect 207140 98590 207360 98640
rect 207140 98520 207150 98590
rect 207350 98520 207360 98590
rect 207140 98480 207360 98520
rect 207140 98410 207150 98480
rect 207350 98410 207360 98480
rect 207140 98360 207360 98410
rect 207640 98590 207860 98640
rect 207640 98520 207650 98590
rect 207850 98520 207860 98590
rect 207640 98480 207860 98520
rect 207640 98410 207650 98480
rect 207850 98410 207860 98480
rect 207640 98360 207860 98410
rect 196000 98350 208000 98360
rect 196000 98150 196020 98350
rect 196090 98150 196410 98350
rect 196480 98150 196520 98350
rect 196590 98150 196910 98350
rect 196980 98150 197020 98350
rect 197090 98150 197410 98350
rect 197480 98150 197520 98350
rect 197590 98150 197910 98350
rect 197980 98150 198020 98350
rect 198090 98150 198410 98350
rect 198480 98150 198520 98350
rect 198590 98150 198910 98350
rect 198980 98150 199020 98350
rect 199090 98150 199410 98350
rect 199480 98150 199520 98350
rect 199590 98150 199910 98350
rect 199980 98150 200020 98350
rect 200090 98150 200410 98350
rect 200480 98150 200520 98350
rect 200590 98150 200910 98350
rect 200980 98150 201020 98350
rect 201090 98150 201410 98350
rect 201480 98150 201520 98350
rect 201590 98150 201910 98350
rect 201980 98150 202020 98350
rect 202090 98150 202410 98350
rect 202480 98150 202520 98350
rect 202590 98150 202910 98350
rect 202980 98150 203020 98350
rect 203090 98150 203410 98350
rect 203480 98150 203520 98350
rect 203590 98150 203910 98350
rect 203980 98150 204020 98350
rect 204090 98150 204410 98350
rect 204480 98150 204520 98350
rect 204590 98150 204910 98350
rect 204980 98150 205020 98350
rect 205090 98150 205410 98350
rect 205480 98150 205520 98350
rect 205590 98150 205910 98350
rect 205980 98150 206020 98350
rect 206090 98150 206410 98350
rect 206480 98150 206520 98350
rect 206590 98150 206910 98350
rect 206980 98150 207020 98350
rect 207090 98150 207410 98350
rect 207480 98150 207520 98350
rect 207590 98150 207910 98350
rect 207980 98150 208000 98350
rect 196000 98140 208000 98150
rect 196140 98090 196360 98140
rect 196140 98020 196150 98090
rect 196350 98020 196360 98090
rect 196140 97980 196360 98020
rect 196140 97910 196150 97980
rect 196350 97910 196360 97980
rect 196140 97860 196360 97910
rect 196640 98090 196860 98140
rect 196640 98020 196650 98090
rect 196850 98020 196860 98090
rect 196640 97980 196860 98020
rect 196640 97910 196650 97980
rect 196850 97910 196860 97980
rect 196640 97860 196860 97910
rect 197140 98090 197360 98140
rect 197140 98020 197150 98090
rect 197350 98020 197360 98090
rect 197140 97980 197360 98020
rect 197140 97910 197150 97980
rect 197350 97910 197360 97980
rect 197140 97860 197360 97910
rect 197640 98090 197860 98140
rect 197640 98020 197650 98090
rect 197850 98020 197860 98090
rect 197640 97980 197860 98020
rect 197640 97910 197650 97980
rect 197850 97910 197860 97980
rect 197640 97860 197860 97910
rect 198140 98090 198360 98140
rect 198140 98020 198150 98090
rect 198350 98020 198360 98090
rect 198140 97980 198360 98020
rect 198140 97910 198150 97980
rect 198350 97910 198360 97980
rect 198140 97860 198360 97910
rect 198640 98090 198860 98140
rect 198640 98020 198650 98090
rect 198850 98020 198860 98090
rect 198640 97980 198860 98020
rect 198640 97910 198650 97980
rect 198850 97910 198860 97980
rect 198640 97860 198860 97910
rect 199140 98090 199360 98140
rect 199140 98020 199150 98090
rect 199350 98020 199360 98090
rect 199140 97980 199360 98020
rect 199140 97910 199150 97980
rect 199350 97910 199360 97980
rect 199140 97860 199360 97910
rect 199640 98090 199860 98140
rect 199640 98020 199650 98090
rect 199850 98020 199860 98090
rect 199640 97980 199860 98020
rect 199640 97910 199650 97980
rect 199850 97910 199860 97980
rect 199640 97860 199860 97910
rect 200140 98090 200360 98140
rect 200140 98020 200150 98090
rect 200350 98020 200360 98090
rect 200140 97980 200360 98020
rect 200140 97910 200150 97980
rect 200350 97910 200360 97980
rect 200140 97860 200360 97910
rect 200640 98090 200860 98140
rect 200640 98020 200650 98090
rect 200850 98020 200860 98090
rect 200640 97980 200860 98020
rect 200640 97910 200650 97980
rect 200850 97910 200860 97980
rect 200640 97860 200860 97910
rect 201140 98090 201360 98140
rect 201140 98020 201150 98090
rect 201350 98020 201360 98090
rect 201140 97980 201360 98020
rect 201140 97910 201150 97980
rect 201350 97910 201360 97980
rect 201140 97860 201360 97910
rect 201640 98090 201860 98140
rect 201640 98020 201650 98090
rect 201850 98020 201860 98090
rect 201640 97980 201860 98020
rect 201640 97910 201650 97980
rect 201850 97910 201860 97980
rect 201640 97860 201860 97910
rect 202140 98090 202360 98140
rect 202140 98020 202150 98090
rect 202350 98020 202360 98090
rect 202140 97980 202360 98020
rect 202140 97910 202150 97980
rect 202350 97910 202360 97980
rect 202140 97860 202360 97910
rect 202640 98090 202860 98140
rect 202640 98020 202650 98090
rect 202850 98020 202860 98090
rect 202640 97980 202860 98020
rect 202640 97910 202650 97980
rect 202850 97910 202860 97980
rect 202640 97860 202860 97910
rect 203140 98090 203360 98140
rect 203140 98020 203150 98090
rect 203350 98020 203360 98090
rect 203140 97980 203360 98020
rect 203140 97910 203150 97980
rect 203350 97910 203360 97980
rect 203140 97860 203360 97910
rect 203640 98090 203860 98140
rect 203640 98020 203650 98090
rect 203850 98020 203860 98090
rect 203640 97980 203860 98020
rect 203640 97910 203650 97980
rect 203850 97910 203860 97980
rect 203640 97860 203860 97910
rect 204140 98090 204360 98140
rect 204140 98020 204150 98090
rect 204350 98020 204360 98090
rect 204140 97980 204360 98020
rect 204140 97910 204150 97980
rect 204350 97910 204360 97980
rect 204140 97860 204360 97910
rect 204640 98090 204860 98140
rect 204640 98020 204650 98090
rect 204850 98020 204860 98090
rect 204640 97980 204860 98020
rect 204640 97910 204650 97980
rect 204850 97910 204860 97980
rect 204640 97860 204860 97910
rect 205140 98090 205360 98140
rect 205140 98020 205150 98090
rect 205350 98020 205360 98090
rect 205140 97980 205360 98020
rect 205140 97910 205150 97980
rect 205350 97910 205360 97980
rect 205140 97860 205360 97910
rect 205640 98090 205860 98140
rect 205640 98020 205650 98090
rect 205850 98020 205860 98090
rect 205640 97980 205860 98020
rect 205640 97910 205650 97980
rect 205850 97910 205860 97980
rect 205640 97860 205860 97910
rect 206140 98090 206360 98140
rect 206140 98020 206150 98090
rect 206350 98020 206360 98090
rect 206140 97980 206360 98020
rect 206140 97910 206150 97980
rect 206350 97910 206360 97980
rect 206140 97860 206360 97910
rect 206640 98090 206860 98140
rect 206640 98020 206650 98090
rect 206850 98020 206860 98090
rect 206640 97980 206860 98020
rect 206640 97910 206650 97980
rect 206850 97910 206860 97980
rect 206640 97860 206860 97910
rect 207140 98090 207360 98140
rect 207140 98020 207150 98090
rect 207350 98020 207360 98090
rect 207140 97980 207360 98020
rect 207140 97910 207150 97980
rect 207350 97910 207360 97980
rect 207140 97860 207360 97910
rect 207640 98090 207860 98140
rect 207640 98020 207650 98090
rect 207850 98020 207860 98090
rect 207640 97980 207860 98020
rect 207640 97910 207650 97980
rect 207850 97910 207860 97980
rect 207640 97860 207860 97910
rect 196000 97850 208000 97860
rect 196000 97650 196020 97850
rect 196090 97650 196410 97850
rect 196480 97650 196520 97850
rect 196590 97650 196910 97850
rect 196980 97650 197020 97850
rect 197090 97650 197410 97850
rect 197480 97650 197520 97850
rect 197590 97650 197910 97850
rect 197980 97650 198020 97850
rect 198090 97650 198410 97850
rect 198480 97650 198520 97850
rect 198590 97650 198910 97850
rect 198980 97650 199020 97850
rect 199090 97650 199410 97850
rect 199480 97650 199520 97850
rect 199590 97650 199910 97850
rect 199980 97650 200020 97850
rect 200090 97650 200410 97850
rect 200480 97650 200520 97850
rect 200590 97650 200910 97850
rect 200980 97650 201020 97850
rect 201090 97650 201410 97850
rect 201480 97650 201520 97850
rect 201590 97650 201910 97850
rect 201980 97650 202020 97850
rect 202090 97650 202410 97850
rect 202480 97650 202520 97850
rect 202590 97650 202910 97850
rect 202980 97650 203020 97850
rect 203090 97650 203410 97850
rect 203480 97650 203520 97850
rect 203590 97650 203910 97850
rect 203980 97650 204020 97850
rect 204090 97650 204410 97850
rect 204480 97650 204520 97850
rect 204590 97650 204910 97850
rect 204980 97650 205020 97850
rect 205090 97650 205410 97850
rect 205480 97650 205520 97850
rect 205590 97650 205910 97850
rect 205980 97650 206020 97850
rect 206090 97650 206410 97850
rect 206480 97650 206520 97850
rect 206590 97650 206910 97850
rect 206980 97650 207020 97850
rect 207090 97650 207410 97850
rect 207480 97650 207520 97850
rect 207590 97650 207910 97850
rect 207980 97650 208000 97850
rect 196000 97640 208000 97650
rect 196140 97590 196360 97640
rect 196140 97520 196150 97590
rect 196350 97520 196360 97590
rect 196140 97480 196360 97520
rect 196140 97410 196150 97480
rect 196350 97410 196360 97480
rect 196140 97360 196360 97410
rect 196640 97590 196860 97640
rect 196640 97520 196650 97590
rect 196850 97520 196860 97590
rect 196640 97480 196860 97520
rect 196640 97410 196650 97480
rect 196850 97410 196860 97480
rect 196640 97360 196860 97410
rect 197140 97590 197360 97640
rect 197140 97520 197150 97590
rect 197350 97520 197360 97590
rect 197140 97480 197360 97520
rect 197140 97410 197150 97480
rect 197350 97410 197360 97480
rect 197140 97360 197360 97410
rect 197640 97590 197860 97640
rect 197640 97520 197650 97590
rect 197850 97520 197860 97590
rect 197640 97480 197860 97520
rect 197640 97410 197650 97480
rect 197850 97410 197860 97480
rect 197640 97360 197860 97410
rect 198140 97590 198360 97640
rect 198140 97520 198150 97590
rect 198350 97520 198360 97590
rect 198140 97480 198360 97520
rect 198140 97410 198150 97480
rect 198350 97410 198360 97480
rect 198140 97360 198360 97410
rect 198640 97590 198860 97640
rect 198640 97520 198650 97590
rect 198850 97520 198860 97590
rect 198640 97480 198860 97520
rect 198640 97410 198650 97480
rect 198850 97410 198860 97480
rect 198640 97360 198860 97410
rect 199140 97590 199360 97640
rect 199140 97520 199150 97590
rect 199350 97520 199360 97590
rect 199140 97480 199360 97520
rect 199140 97410 199150 97480
rect 199350 97410 199360 97480
rect 199140 97360 199360 97410
rect 199640 97590 199860 97640
rect 199640 97520 199650 97590
rect 199850 97520 199860 97590
rect 199640 97480 199860 97520
rect 199640 97410 199650 97480
rect 199850 97410 199860 97480
rect 199640 97360 199860 97410
rect 200140 97590 200360 97640
rect 200140 97520 200150 97590
rect 200350 97520 200360 97590
rect 200140 97480 200360 97520
rect 200140 97410 200150 97480
rect 200350 97410 200360 97480
rect 200140 97360 200360 97410
rect 200640 97590 200860 97640
rect 200640 97520 200650 97590
rect 200850 97520 200860 97590
rect 200640 97480 200860 97520
rect 200640 97410 200650 97480
rect 200850 97410 200860 97480
rect 200640 97360 200860 97410
rect 201140 97590 201360 97640
rect 201140 97520 201150 97590
rect 201350 97520 201360 97590
rect 201140 97480 201360 97520
rect 201140 97410 201150 97480
rect 201350 97410 201360 97480
rect 201140 97360 201360 97410
rect 201640 97590 201860 97640
rect 201640 97520 201650 97590
rect 201850 97520 201860 97590
rect 201640 97480 201860 97520
rect 201640 97410 201650 97480
rect 201850 97410 201860 97480
rect 201640 97360 201860 97410
rect 202140 97590 202360 97640
rect 202140 97520 202150 97590
rect 202350 97520 202360 97590
rect 202140 97480 202360 97520
rect 202140 97410 202150 97480
rect 202350 97410 202360 97480
rect 202140 97360 202360 97410
rect 202640 97590 202860 97640
rect 202640 97520 202650 97590
rect 202850 97520 202860 97590
rect 202640 97480 202860 97520
rect 202640 97410 202650 97480
rect 202850 97410 202860 97480
rect 202640 97360 202860 97410
rect 203140 97590 203360 97640
rect 203140 97520 203150 97590
rect 203350 97520 203360 97590
rect 203140 97480 203360 97520
rect 203140 97410 203150 97480
rect 203350 97410 203360 97480
rect 203140 97360 203360 97410
rect 203640 97590 203860 97640
rect 203640 97520 203650 97590
rect 203850 97520 203860 97590
rect 203640 97480 203860 97520
rect 203640 97410 203650 97480
rect 203850 97410 203860 97480
rect 203640 97360 203860 97410
rect 204140 97590 204360 97640
rect 204140 97520 204150 97590
rect 204350 97520 204360 97590
rect 204140 97480 204360 97520
rect 204140 97410 204150 97480
rect 204350 97410 204360 97480
rect 204140 97360 204360 97410
rect 204640 97590 204860 97640
rect 204640 97520 204650 97590
rect 204850 97520 204860 97590
rect 204640 97480 204860 97520
rect 204640 97410 204650 97480
rect 204850 97410 204860 97480
rect 204640 97360 204860 97410
rect 205140 97590 205360 97640
rect 205140 97520 205150 97590
rect 205350 97520 205360 97590
rect 205140 97480 205360 97520
rect 205140 97410 205150 97480
rect 205350 97410 205360 97480
rect 205140 97360 205360 97410
rect 205640 97590 205860 97640
rect 205640 97520 205650 97590
rect 205850 97520 205860 97590
rect 205640 97480 205860 97520
rect 205640 97410 205650 97480
rect 205850 97410 205860 97480
rect 205640 97360 205860 97410
rect 206140 97590 206360 97640
rect 206140 97520 206150 97590
rect 206350 97520 206360 97590
rect 206140 97480 206360 97520
rect 206140 97410 206150 97480
rect 206350 97410 206360 97480
rect 206140 97360 206360 97410
rect 206640 97590 206860 97640
rect 206640 97520 206650 97590
rect 206850 97520 206860 97590
rect 206640 97480 206860 97520
rect 206640 97410 206650 97480
rect 206850 97410 206860 97480
rect 206640 97360 206860 97410
rect 207140 97590 207360 97640
rect 207140 97520 207150 97590
rect 207350 97520 207360 97590
rect 207140 97480 207360 97520
rect 207140 97410 207150 97480
rect 207350 97410 207360 97480
rect 207140 97360 207360 97410
rect 207640 97590 207860 97640
rect 207640 97520 207650 97590
rect 207850 97520 207860 97590
rect 207640 97480 207860 97520
rect 207640 97410 207650 97480
rect 207850 97410 207860 97480
rect 207640 97360 207860 97410
rect 196000 97350 208000 97360
rect 196000 97150 196020 97350
rect 196090 97150 196410 97350
rect 196480 97150 196520 97350
rect 196590 97150 196910 97350
rect 196980 97150 197020 97350
rect 197090 97150 197410 97350
rect 197480 97150 197520 97350
rect 197590 97150 197910 97350
rect 197980 97150 198020 97350
rect 198090 97150 198410 97350
rect 198480 97150 198520 97350
rect 198590 97150 198910 97350
rect 198980 97150 199020 97350
rect 199090 97150 199410 97350
rect 199480 97150 199520 97350
rect 199590 97150 199910 97350
rect 199980 97150 200020 97350
rect 200090 97150 200410 97350
rect 200480 97150 200520 97350
rect 200590 97150 200910 97350
rect 200980 97150 201020 97350
rect 201090 97150 201410 97350
rect 201480 97150 201520 97350
rect 201590 97150 201910 97350
rect 201980 97150 202020 97350
rect 202090 97150 202410 97350
rect 202480 97150 202520 97350
rect 202590 97150 202910 97350
rect 202980 97150 203020 97350
rect 203090 97150 203410 97350
rect 203480 97150 203520 97350
rect 203590 97150 203910 97350
rect 203980 97150 204020 97350
rect 204090 97150 204410 97350
rect 204480 97150 204520 97350
rect 204590 97150 204910 97350
rect 204980 97150 205020 97350
rect 205090 97150 205410 97350
rect 205480 97150 205520 97350
rect 205590 97150 205910 97350
rect 205980 97150 206020 97350
rect 206090 97150 206410 97350
rect 206480 97150 206520 97350
rect 206590 97150 206910 97350
rect 206980 97150 207020 97350
rect 207090 97150 207410 97350
rect 207480 97150 207520 97350
rect 207590 97150 207910 97350
rect 207980 97150 208000 97350
rect 196000 97140 208000 97150
rect 196140 97090 196360 97140
rect 196140 97020 196150 97090
rect 196350 97020 196360 97090
rect 196140 96980 196360 97020
rect 196140 96910 196150 96980
rect 196350 96910 196360 96980
rect 196140 96860 196360 96910
rect 196640 97090 196860 97140
rect 196640 97020 196650 97090
rect 196850 97020 196860 97090
rect 196640 96980 196860 97020
rect 196640 96910 196650 96980
rect 196850 96910 196860 96980
rect 196640 96860 196860 96910
rect 197140 97090 197360 97140
rect 197140 97020 197150 97090
rect 197350 97020 197360 97090
rect 197140 96980 197360 97020
rect 197140 96910 197150 96980
rect 197350 96910 197360 96980
rect 197140 96860 197360 96910
rect 197640 97090 197860 97140
rect 197640 97020 197650 97090
rect 197850 97020 197860 97090
rect 197640 96980 197860 97020
rect 197640 96910 197650 96980
rect 197850 96910 197860 96980
rect 197640 96860 197860 96910
rect 198140 97090 198360 97140
rect 198140 97020 198150 97090
rect 198350 97020 198360 97090
rect 198140 96980 198360 97020
rect 198140 96910 198150 96980
rect 198350 96910 198360 96980
rect 198140 96860 198360 96910
rect 198640 97090 198860 97140
rect 198640 97020 198650 97090
rect 198850 97020 198860 97090
rect 198640 96980 198860 97020
rect 198640 96910 198650 96980
rect 198850 96910 198860 96980
rect 198640 96860 198860 96910
rect 199140 97090 199360 97140
rect 199140 97020 199150 97090
rect 199350 97020 199360 97090
rect 199140 96980 199360 97020
rect 199140 96910 199150 96980
rect 199350 96910 199360 96980
rect 199140 96860 199360 96910
rect 199640 97090 199860 97140
rect 199640 97020 199650 97090
rect 199850 97020 199860 97090
rect 199640 96980 199860 97020
rect 199640 96910 199650 96980
rect 199850 96910 199860 96980
rect 199640 96860 199860 96910
rect 200140 97090 200360 97140
rect 200140 97020 200150 97090
rect 200350 97020 200360 97090
rect 200140 96980 200360 97020
rect 200140 96910 200150 96980
rect 200350 96910 200360 96980
rect 200140 96860 200360 96910
rect 200640 97090 200860 97140
rect 200640 97020 200650 97090
rect 200850 97020 200860 97090
rect 200640 96980 200860 97020
rect 200640 96910 200650 96980
rect 200850 96910 200860 96980
rect 200640 96860 200860 96910
rect 201140 97090 201360 97140
rect 201140 97020 201150 97090
rect 201350 97020 201360 97090
rect 201140 96980 201360 97020
rect 201140 96910 201150 96980
rect 201350 96910 201360 96980
rect 201140 96860 201360 96910
rect 201640 97090 201860 97140
rect 201640 97020 201650 97090
rect 201850 97020 201860 97090
rect 201640 96980 201860 97020
rect 201640 96910 201650 96980
rect 201850 96910 201860 96980
rect 201640 96860 201860 96910
rect 202140 97090 202360 97140
rect 202140 97020 202150 97090
rect 202350 97020 202360 97090
rect 202140 96980 202360 97020
rect 202140 96910 202150 96980
rect 202350 96910 202360 96980
rect 202140 96860 202360 96910
rect 202640 97090 202860 97140
rect 202640 97020 202650 97090
rect 202850 97020 202860 97090
rect 202640 96980 202860 97020
rect 202640 96910 202650 96980
rect 202850 96910 202860 96980
rect 202640 96860 202860 96910
rect 203140 97090 203360 97140
rect 203140 97020 203150 97090
rect 203350 97020 203360 97090
rect 203140 96980 203360 97020
rect 203140 96910 203150 96980
rect 203350 96910 203360 96980
rect 203140 96860 203360 96910
rect 203640 97090 203860 97140
rect 203640 97020 203650 97090
rect 203850 97020 203860 97090
rect 203640 96980 203860 97020
rect 203640 96910 203650 96980
rect 203850 96910 203860 96980
rect 203640 96860 203860 96910
rect 204140 97090 204360 97140
rect 204140 97020 204150 97090
rect 204350 97020 204360 97090
rect 204140 96980 204360 97020
rect 204140 96910 204150 96980
rect 204350 96910 204360 96980
rect 204140 96860 204360 96910
rect 204640 97090 204860 97140
rect 204640 97020 204650 97090
rect 204850 97020 204860 97090
rect 204640 96980 204860 97020
rect 204640 96910 204650 96980
rect 204850 96910 204860 96980
rect 204640 96860 204860 96910
rect 205140 97090 205360 97140
rect 205140 97020 205150 97090
rect 205350 97020 205360 97090
rect 205140 96980 205360 97020
rect 205140 96910 205150 96980
rect 205350 96910 205360 96980
rect 205140 96860 205360 96910
rect 205640 97090 205860 97140
rect 205640 97020 205650 97090
rect 205850 97020 205860 97090
rect 205640 96980 205860 97020
rect 205640 96910 205650 96980
rect 205850 96910 205860 96980
rect 205640 96860 205860 96910
rect 206140 97090 206360 97140
rect 206140 97020 206150 97090
rect 206350 97020 206360 97090
rect 206140 96980 206360 97020
rect 206140 96910 206150 96980
rect 206350 96910 206360 96980
rect 206140 96860 206360 96910
rect 206640 97090 206860 97140
rect 206640 97020 206650 97090
rect 206850 97020 206860 97090
rect 206640 96980 206860 97020
rect 206640 96910 206650 96980
rect 206850 96910 206860 96980
rect 206640 96860 206860 96910
rect 207140 97090 207360 97140
rect 207140 97020 207150 97090
rect 207350 97020 207360 97090
rect 207140 96980 207360 97020
rect 207140 96910 207150 96980
rect 207350 96910 207360 96980
rect 207140 96860 207360 96910
rect 207640 97090 207860 97140
rect 207640 97020 207650 97090
rect 207850 97020 207860 97090
rect 207640 96980 207860 97020
rect 207640 96910 207650 96980
rect 207850 96910 207860 96980
rect 207640 96860 207860 96910
rect 196000 96850 208000 96860
rect 196000 96650 196020 96850
rect 196090 96650 196410 96850
rect 196480 96650 196520 96850
rect 196590 96650 196910 96850
rect 196980 96650 197020 96850
rect 197090 96650 197410 96850
rect 197480 96650 197520 96850
rect 197590 96650 197910 96850
rect 197980 96650 198020 96850
rect 198090 96650 198410 96850
rect 198480 96650 198520 96850
rect 198590 96650 198910 96850
rect 198980 96650 199020 96850
rect 199090 96650 199410 96850
rect 199480 96650 199520 96850
rect 199590 96650 199910 96850
rect 199980 96650 200020 96850
rect 200090 96650 200410 96850
rect 200480 96650 200520 96850
rect 200590 96650 200910 96850
rect 200980 96650 201020 96850
rect 201090 96650 201410 96850
rect 201480 96650 201520 96850
rect 201590 96650 201910 96850
rect 201980 96650 202020 96850
rect 202090 96650 202410 96850
rect 202480 96650 202520 96850
rect 202590 96650 202910 96850
rect 202980 96650 203020 96850
rect 203090 96650 203410 96850
rect 203480 96650 203520 96850
rect 203590 96650 203910 96850
rect 203980 96650 204020 96850
rect 204090 96650 204410 96850
rect 204480 96650 204520 96850
rect 204590 96650 204910 96850
rect 204980 96650 205020 96850
rect 205090 96650 205410 96850
rect 205480 96650 205520 96850
rect 205590 96650 205910 96850
rect 205980 96650 206020 96850
rect 206090 96650 206410 96850
rect 206480 96650 206520 96850
rect 206590 96650 206910 96850
rect 206980 96650 207020 96850
rect 207090 96650 207410 96850
rect 207480 96650 207520 96850
rect 207590 96650 207910 96850
rect 207980 96650 208000 96850
rect 196000 96640 208000 96650
rect 196140 96590 196360 96640
rect 196140 96520 196150 96590
rect 196350 96520 196360 96590
rect 196140 96480 196360 96520
rect 196140 96410 196150 96480
rect 196350 96410 196360 96480
rect 196140 96360 196360 96410
rect 196640 96590 196860 96640
rect 196640 96520 196650 96590
rect 196850 96520 196860 96590
rect 196640 96480 196860 96520
rect 196640 96410 196650 96480
rect 196850 96410 196860 96480
rect 196640 96360 196860 96410
rect 197140 96590 197360 96640
rect 197140 96520 197150 96590
rect 197350 96520 197360 96590
rect 197140 96480 197360 96520
rect 197140 96410 197150 96480
rect 197350 96410 197360 96480
rect 197140 96360 197360 96410
rect 197640 96590 197860 96640
rect 197640 96520 197650 96590
rect 197850 96520 197860 96590
rect 197640 96480 197860 96520
rect 197640 96410 197650 96480
rect 197850 96410 197860 96480
rect 197640 96360 197860 96410
rect 198140 96590 198360 96640
rect 198140 96520 198150 96590
rect 198350 96520 198360 96590
rect 198140 96480 198360 96520
rect 198140 96410 198150 96480
rect 198350 96410 198360 96480
rect 198140 96360 198360 96410
rect 198640 96590 198860 96640
rect 198640 96520 198650 96590
rect 198850 96520 198860 96590
rect 198640 96480 198860 96520
rect 198640 96410 198650 96480
rect 198850 96410 198860 96480
rect 198640 96360 198860 96410
rect 199140 96590 199360 96640
rect 199140 96520 199150 96590
rect 199350 96520 199360 96590
rect 199140 96480 199360 96520
rect 199140 96410 199150 96480
rect 199350 96410 199360 96480
rect 199140 96360 199360 96410
rect 199640 96590 199860 96640
rect 199640 96520 199650 96590
rect 199850 96520 199860 96590
rect 199640 96480 199860 96520
rect 199640 96410 199650 96480
rect 199850 96410 199860 96480
rect 199640 96360 199860 96410
rect 200140 96590 200360 96640
rect 200140 96520 200150 96590
rect 200350 96520 200360 96590
rect 200140 96480 200360 96520
rect 200140 96410 200150 96480
rect 200350 96410 200360 96480
rect 200140 96360 200360 96410
rect 200640 96590 200860 96640
rect 200640 96520 200650 96590
rect 200850 96520 200860 96590
rect 200640 96480 200860 96520
rect 200640 96410 200650 96480
rect 200850 96410 200860 96480
rect 200640 96360 200860 96410
rect 201140 96590 201360 96640
rect 201140 96520 201150 96590
rect 201350 96520 201360 96590
rect 201140 96480 201360 96520
rect 201140 96410 201150 96480
rect 201350 96410 201360 96480
rect 201140 96360 201360 96410
rect 201640 96590 201860 96640
rect 201640 96520 201650 96590
rect 201850 96520 201860 96590
rect 201640 96480 201860 96520
rect 201640 96410 201650 96480
rect 201850 96410 201860 96480
rect 201640 96360 201860 96410
rect 202140 96590 202360 96640
rect 202140 96520 202150 96590
rect 202350 96520 202360 96590
rect 202140 96480 202360 96520
rect 202140 96410 202150 96480
rect 202350 96410 202360 96480
rect 202140 96360 202360 96410
rect 202640 96590 202860 96640
rect 202640 96520 202650 96590
rect 202850 96520 202860 96590
rect 202640 96480 202860 96520
rect 202640 96410 202650 96480
rect 202850 96410 202860 96480
rect 202640 96360 202860 96410
rect 203140 96590 203360 96640
rect 203140 96520 203150 96590
rect 203350 96520 203360 96590
rect 203140 96480 203360 96520
rect 203140 96410 203150 96480
rect 203350 96410 203360 96480
rect 203140 96360 203360 96410
rect 203640 96590 203860 96640
rect 203640 96520 203650 96590
rect 203850 96520 203860 96590
rect 203640 96480 203860 96520
rect 203640 96410 203650 96480
rect 203850 96410 203860 96480
rect 203640 96360 203860 96410
rect 204140 96590 204360 96640
rect 204140 96520 204150 96590
rect 204350 96520 204360 96590
rect 204140 96480 204360 96520
rect 204140 96410 204150 96480
rect 204350 96410 204360 96480
rect 204140 96360 204360 96410
rect 204640 96590 204860 96640
rect 204640 96520 204650 96590
rect 204850 96520 204860 96590
rect 204640 96480 204860 96520
rect 204640 96410 204650 96480
rect 204850 96410 204860 96480
rect 204640 96360 204860 96410
rect 205140 96590 205360 96640
rect 205140 96520 205150 96590
rect 205350 96520 205360 96590
rect 205140 96480 205360 96520
rect 205140 96410 205150 96480
rect 205350 96410 205360 96480
rect 205140 96360 205360 96410
rect 205640 96590 205860 96640
rect 205640 96520 205650 96590
rect 205850 96520 205860 96590
rect 205640 96480 205860 96520
rect 205640 96410 205650 96480
rect 205850 96410 205860 96480
rect 205640 96360 205860 96410
rect 206140 96590 206360 96640
rect 206140 96520 206150 96590
rect 206350 96520 206360 96590
rect 206140 96480 206360 96520
rect 206140 96410 206150 96480
rect 206350 96410 206360 96480
rect 206140 96360 206360 96410
rect 206640 96590 206860 96640
rect 206640 96520 206650 96590
rect 206850 96520 206860 96590
rect 206640 96480 206860 96520
rect 206640 96410 206650 96480
rect 206850 96410 206860 96480
rect 206640 96360 206860 96410
rect 207140 96590 207360 96640
rect 207140 96520 207150 96590
rect 207350 96520 207360 96590
rect 207140 96480 207360 96520
rect 207140 96410 207150 96480
rect 207350 96410 207360 96480
rect 207140 96360 207360 96410
rect 207640 96590 207860 96640
rect 207640 96520 207650 96590
rect 207850 96520 207860 96590
rect 207640 96480 207860 96520
rect 207640 96410 207650 96480
rect 207850 96410 207860 96480
rect 207640 96360 207860 96410
rect 196000 96350 208000 96360
rect 196000 96150 196020 96350
rect 196090 96150 196410 96350
rect 196480 96150 196520 96350
rect 196590 96150 196910 96350
rect 196980 96150 197020 96350
rect 197090 96150 197410 96350
rect 197480 96150 197520 96350
rect 197590 96150 197910 96350
rect 197980 96150 198020 96350
rect 198090 96150 198410 96350
rect 198480 96150 198520 96350
rect 198590 96150 198910 96350
rect 198980 96150 199020 96350
rect 199090 96150 199410 96350
rect 199480 96150 199520 96350
rect 199590 96150 199910 96350
rect 199980 96150 200020 96350
rect 200090 96150 200410 96350
rect 200480 96150 200520 96350
rect 200590 96150 200910 96350
rect 200980 96150 201020 96350
rect 201090 96150 201410 96350
rect 201480 96150 201520 96350
rect 201590 96150 201910 96350
rect 201980 96150 202020 96350
rect 202090 96150 202410 96350
rect 202480 96150 202520 96350
rect 202590 96150 202910 96350
rect 202980 96150 203020 96350
rect 203090 96150 203410 96350
rect 203480 96150 203520 96350
rect 203590 96150 203910 96350
rect 203980 96150 204020 96350
rect 204090 96150 204410 96350
rect 204480 96150 204520 96350
rect 204590 96150 204910 96350
rect 204980 96150 205020 96350
rect 205090 96150 205410 96350
rect 205480 96150 205520 96350
rect 205590 96150 205910 96350
rect 205980 96150 206020 96350
rect 206090 96150 206410 96350
rect 206480 96150 206520 96350
rect 206590 96150 206910 96350
rect 206980 96150 207020 96350
rect 207090 96150 207410 96350
rect 207480 96150 207520 96350
rect 207590 96150 207910 96350
rect 207980 96150 208000 96350
rect 196000 96140 208000 96150
rect 196140 96090 196360 96140
rect 196140 96020 196150 96090
rect 196350 96020 196360 96090
rect 196140 95980 196360 96020
rect 196140 95910 196150 95980
rect 196350 95910 196360 95980
rect 196140 95860 196360 95910
rect 196640 96090 196860 96140
rect 196640 96020 196650 96090
rect 196850 96020 196860 96090
rect 196640 95980 196860 96020
rect 196640 95910 196650 95980
rect 196850 95910 196860 95980
rect 196640 95860 196860 95910
rect 197140 96090 197360 96140
rect 197140 96020 197150 96090
rect 197350 96020 197360 96090
rect 197140 95980 197360 96020
rect 197140 95910 197150 95980
rect 197350 95910 197360 95980
rect 197140 95860 197360 95910
rect 197640 96090 197860 96140
rect 197640 96020 197650 96090
rect 197850 96020 197860 96090
rect 197640 95980 197860 96020
rect 197640 95910 197650 95980
rect 197850 95910 197860 95980
rect 197640 95860 197860 95910
rect 198140 96090 198360 96140
rect 198140 96020 198150 96090
rect 198350 96020 198360 96090
rect 198140 95980 198360 96020
rect 198140 95910 198150 95980
rect 198350 95910 198360 95980
rect 198140 95860 198360 95910
rect 198640 96090 198860 96140
rect 198640 96020 198650 96090
rect 198850 96020 198860 96090
rect 198640 95980 198860 96020
rect 198640 95910 198650 95980
rect 198850 95910 198860 95980
rect 198640 95860 198860 95910
rect 199140 96090 199360 96140
rect 199140 96020 199150 96090
rect 199350 96020 199360 96090
rect 199140 95980 199360 96020
rect 199140 95910 199150 95980
rect 199350 95910 199360 95980
rect 199140 95860 199360 95910
rect 199640 96090 199860 96140
rect 199640 96020 199650 96090
rect 199850 96020 199860 96090
rect 199640 95980 199860 96020
rect 199640 95910 199650 95980
rect 199850 95910 199860 95980
rect 199640 95860 199860 95910
rect 200140 96090 200360 96140
rect 200140 96020 200150 96090
rect 200350 96020 200360 96090
rect 200140 95980 200360 96020
rect 200140 95910 200150 95980
rect 200350 95910 200360 95980
rect 200140 95860 200360 95910
rect 200640 96090 200860 96140
rect 200640 96020 200650 96090
rect 200850 96020 200860 96090
rect 200640 95980 200860 96020
rect 200640 95910 200650 95980
rect 200850 95910 200860 95980
rect 200640 95860 200860 95910
rect 201140 96090 201360 96140
rect 201140 96020 201150 96090
rect 201350 96020 201360 96090
rect 201140 95980 201360 96020
rect 201140 95910 201150 95980
rect 201350 95910 201360 95980
rect 201140 95860 201360 95910
rect 201640 96090 201860 96140
rect 201640 96020 201650 96090
rect 201850 96020 201860 96090
rect 201640 95980 201860 96020
rect 201640 95910 201650 95980
rect 201850 95910 201860 95980
rect 201640 95860 201860 95910
rect 202140 96090 202360 96140
rect 202140 96020 202150 96090
rect 202350 96020 202360 96090
rect 202140 95980 202360 96020
rect 202140 95910 202150 95980
rect 202350 95910 202360 95980
rect 202140 95860 202360 95910
rect 202640 96090 202860 96140
rect 202640 96020 202650 96090
rect 202850 96020 202860 96090
rect 202640 95980 202860 96020
rect 202640 95910 202650 95980
rect 202850 95910 202860 95980
rect 202640 95860 202860 95910
rect 203140 96090 203360 96140
rect 203140 96020 203150 96090
rect 203350 96020 203360 96090
rect 203140 95980 203360 96020
rect 203140 95910 203150 95980
rect 203350 95910 203360 95980
rect 203140 95860 203360 95910
rect 203640 96090 203860 96140
rect 203640 96020 203650 96090
rect 203850 96020 203860 96090
rect 203640 95980 203860 96020
rect 203640 95910 203650 95980
rect 203850 95910 203860 95980
rect 203640 95860 203860 95910
rect 204140 96090 204360 96140
rect 204140 96020 204150 96090
rect 204350 96020 204360 96090
rect 204140 95980 204360 96020
rect 204140 95910 204150 95980
rect 204350 95910 204360 95980
rect 204140 95860 204360 95910
rect 204640 96090 204860 96140
rect 204640 96020 204650 96090
rect 204850 96020 204860 96090
rect 204640 95980 204860 96020
rect 204640 95910 204650 95980
rect 204850 95910 204860 95980
rect 204640 95860 204860 95910
rect 205140 96090 205360 96140
rect 205140 96020 205150 96090
rect 205350 96020 205360 96090
rect 205140 95980 205360 96020
rect 205140 95910 205150 95980
rect 205350 95910 205360 95980
rect 205140 95860 205360 95910
rect 205640 96090 205860 96140
rect 205640 96020 205650 96090
rect 205850 96020 205860 96090
rect 205640 95980 205860 96020
rect 205640 95910 205650 95980
rect 205850 95910 205860 95980
rect 205640 95860 205860 95910
rect 206140 96090 206360 96140
rect 206140 96020 206150 96090
rect 206350 96020 206360 96090
rect 206140 95980 206360 96020
rect 206140 95910 206150 95980
rect 206350 95910 206360 95980
rect 206140 95860 206360 95910
rect 206640 96090 206860 96140
rect 206640 96020 206650 96090
rect 206850 96020 206860 96090
rect 206640 95980 206860 96020
rect 206640 95910 206650 95980
rect 206850 95910 206860 95980
rect 206640 95860 206860 95910
rect 207140 96090 207360 96140
rect 207140 96020 207150 96090
rect 207350 96020 207360 96090
rect 207140 95980 207360 96020
rect 207140 95910 207150 95980
rect 207350 95910 207360 95980
rect 207140 95860 207360 95910
rect 207640 96090 207860 96140
rect 207640 96020 207650 96090
rect 207850 96020 207860 96090
rect 207640 95980 207860 96020
rect 207640 95910 207650 95980
rect 207850 95910 207860 95980
rect 207640 95860 207860 95910
rect 196000 95850 208000 95860
rect 196000 95650 196020 95850
rect 196090 95650 196410 95850
rect 196480 95650 196520 95850
rect 196590 95650 196910 95850
rect 196980 95650 197020 95850
rect 197090 95650 197410 95850
rect 197480 95650 197520 95850
rect 197590 95650 197910 95850
rect 197980 95650 198020 95850
rect 198090 95650 198410 95850
rect 198480 95650 198520 95850
rect 198590 95650 198910 95850
rect 198980 95650 199020 95850
rect 199090 95650 199410 95850
rect 199480 95650 199520 95850
rect 199590 95650 199910 95850
rect 199980 95650 200020 95850
rect 200090 95650 200410 95850
rect 200480 95650 200520 95850
rect 200590 95650 200910 95850
rect 200980 95650 201020 95850
rect 201090 95650 201410 95850
rect 201480 95650 201520 95850
rect 201590 95650 201910 95850
rect 201980 95650 202020 95850
rect 202090 95650 202410 95850
rect 202480 95650 202520 95850
rect 202590 95650 202910 95850
rect 202980 95650 203020 95850
rect 203090 95650 203410 95850
rect 203480 95650 203520 95850
rect 203590 95650 203910 95850
rect 203980 95650 204020 95850
rect 204090 95650 204410 95850
rect 204480 95650 204520 95850
rect 204590 95650 204910 95850
rect 204980 95650 205020 95850
rect 205090 95650 205410 95850
rect 205480 95650 205520 95850
rect 205590 95650 205910 95850
rect 205980 95650 206020 95850
rect 206090 95650 206410 95850
rect 206480 95650 206520 95850
rect 206590 95650 206910 95850
rect 206980 95650 207020 95850
rect 207090 95650 207410 95850
rect 207480 95650 207520 95850
rect 207590 95650 207910 95850
rect 207980 95650 208000 95850
rect 196000 95640 208000 95650
rect 196140 95590 196360 95640
rect 196140 95520 196150 95590
rect 196350 95520 196360 95590
rect 196140 95480 196360 95520
rect 196140 95410 196150 95480
rect 196350 95410 196360 95480
rect 196140 95360 196360 95410
rect 196640 95590 196860 95640
rect 196640 95520 196650 95590
rect 196850 95520 196860 95590
rect 196640 95480 196860 95520
rect 196640 95410 196650 95480
rect 196850 95410 196860 95480
rect 196640 95360 196860 95410
rect 197140 95590 197360 95640
rect 197140 95520 197150 95590
rect 197350 95520 197360 95590
rect 197140 95480 197360 95520
rect 197140 95410 197150 95480
rect 197350 95410 197360 95480
rect 197140 95360 197360 95410
rect 197640 95590 197860 95640
rect 197640 95520 197650 95590
rect 197850 95520 197860 95590
rect 197640 95480 197860 95520
rect 197640 95410 197650 95480
rect 197850 95410 197860 95480
rect 197640 95360 197860 95410
rect 198140 95590 198360 95640
rect 198140 95520 198150 95590
rect 198350 95520 198360 95590
rect 198140 95480 198360 95520
rect 198140 95410 198150 95480
rect 198350 95410 198360 95480
rect 198140 95360 198360 95410
rect 198640 95590 198860 95640
rect 198640 95520 198650 95590
rect 198850 95520 198860 95590
rect 198640 95480 198860 95520
rect 198640 95410 198650 95480
rect 198850 95410 198860 95480
rect 198640 95360 198860 95410
rect 199140 95590 199360 95640
rect 199140 95520 199150 95590
rect 199350 95520 199360 95590
rect 199140 95480 199360 95520
rect 199140 95410 199150 95480
rect 199350 95410 199360 95480
rect 199140 95360 199360 95410
rect 199640 95590 199860 95640
rect 199640 95520 199650 95590
rect 199850 95520 199860 95590
rect 199640 95480 199860 95520
rect 199640 95410 199650 95480
rect 199850 95410 199860 95480
rect 199640 95360 199860 95410
rect 200140 95590 200360 95640
rect 200140 95520 200150 95590
rect 200350 95520 200360 95590
rect 200140 95480 200360 95520
rect 200140 95410 200150 95480
rect 200350 95410 200360 95480
rect 200140 95360 200360 95410
rect 200640 95590 200860 95640
rect 200640 95520 200650 95590
rect 200850 95520 200860 95590
rect 200640 95480 200860 95520
rect 200640 95410 200650 95480
rect 200850 95410 200860 95480
rect 200640 95360 200860 95410
rect 201140 95590 201360 95640
rect 201140 95520 201150 95590
rect 201350 95520 201360 95590
rect 201140 95480 201360 95520
rect 201140 95410 201150 95480
rect 201350 95410 201360 95480
rect 201140 95360 201360 95410
rect 201640 95590 201860 95640
rect 201640 95520 201650 95590
rect 201850 95520 201860 95590
rect 201640 95480 201860 95520
rect 201640 95410 201650 95480
rect 201850 95410 201860 95480
rect 201640 95360 201860 95410
rect 202140 95590 202360 95640
rect 202140 95520 202150 95590
rect 202350 95520 202360 95590
rect 202140 95480 202360 95520
rect 202140 95410 202150 95480
rect 202350 95410 202360 95480
rect 202140 95360 202360 95410
rect 202640 95590 202860 95640
rect 202640 95520 202650 95590
rect 202850 95520 202860 95590
rect 202640 95480 202860 95520
rect 202640 95410 202650 95480
rect 202850 95410 202860 95480
rect 202640 95360 202860 95410
rect 203140 95590 203360 95640
rect 203140 95520 203150 95590
rect 203350 95520 203360 95590
rect 203140 95480 203360 95520
rect 203140 95410 203150 95480
rect 203350 95410 203360 95480
rect 203140 95360 203360 95410
rect 203640 95590 203860 95640
rect 203640 95520 203650 95590
rect 203850 95520 203860 95590
rect 203640 95480 203860 95520
rect 203640 95410 203650 95480
rect 203850 95410 203860 95480
rect 203640 95360 203860 95410
rect 204140 95590 204360 95640
rect 204140 95520 204150 95590
rect 204350 95520 204360 95590
rect 204140 95480 204360 95520
rect 204140 95410 204150 95480
rect 204350 95410 204360 95480
rect 204140 95360 204360 95410
rect 204640 95590 204860 95640
rect 204640 95520 204650 95590
rect 204850 95520 204860 95590
rect 204640 95480 204860 95520
rect 204640 95410 204650 95480
rect 204850 95410 204860 95480
rect 204640 95360 204860 95410
rect 205140 95590 205360 95640
rect 205140 95520 205150 95590
rect 205350 95520 205360 95590
rect 205140 95480 205360 95520
rect 205140 95410 205150 95480
rect 205350 95410 205360 95480
rect 205140 95360 205360 95410
rect 205640 95590 205860 95640
rect 205640 95520 205650 95590
rect 205850 95520 205860 95590
rect 205640 95480 205860 95520
rect 205640 95410 205650 95480
rect 205850 95410 205860 95480
rect 205640 95360 205860 95410
rect 206140 95590 206360 95640
rect 206140 95520 206150 95590
rect 206350 95520 206360 95590
rect 206140 95480 206360 95520
rect 206140 95410 206150 95480
rect 206350 95410 206360 95480
rect 206140 95360 206360 95410
rect 206640 95590 206860 95640
rect 206640 95520 206650 95590
rect 206850 95520 206860 95590
rect 206640 95480 206860 95520
rect 206640 95410 206650 95480
rect 206850 95410 206860 95480
rect 206640 95360 206860 95410
rect 207140 95590 207360 95640
rect 207140 95520 207150 95590
rect 207350 95520 207360 95590
rect 207140 95480 207360 95520
rect 207140 95410 207150 95480
rect 207350 95410 207360 95480
rect 207140 95360 207360 95410
rect 207640 95590 207860 95640
rect 207640 95520 207650 95590
rect 207850 95520 207860 95590
rect 207640 95480 207860 95520
rect 207640 95410 207650 95480
rect 207850 95410 207860 95480
rect 207640 95360 207860 95410
rect 196000 95350 208000 95360
rect 196000 95150 196020 95350
rect 196090 95150 196410 95350
rect 196480 95150 196520 95350
rect 196590 95150 196910 95350
rect 196980 95150 197020 95350
rect 197090 95150 197410 95350
rect 197480 95150 197520 95350
rect 197590 95150 197910 95350
rect 197980 95150 198020 95350
rect 198090 95150 198410 95350
rect 198480 95150 198520 95350
rect 198590 95150 198910 95350
rect 198980 95150 199020 95350
rect 199090 95150 199410 95350
rect 199480 95150 199520 95350
rect 199590 95150 199910 95350
rect 199980 95150 200020 95350
rect 200090 95150 200410 95350
rect 200480 95150 200520 95350
rect 200590 95150 200910 95350
rect 200980 95150 201020 95350
rect 201090 95150 201410 95350
rect 201480 95150 201520 95350
rect 201590 95150 201910 95350
rect 201980 95150 202020 95350
rect 202090 95150 202410 95350
rect 202480 95150 202520 95350
rect 202590 95150 202910 95350
rect 202980 95150 203020 95350
rect 203090 95150 203410 95350
rect 203480 95150 203520 95350
rect 203590 95150 203910 95350
rect 203980 95150 204020 95350
rect 204090 95150 204410 95350
rect 204480 95150 204520 95350
rect 204590 95150 204910 95350
rect 204980 95150 205020 95350
rect 205090 95150 205410 95350
rect 205480 95150 205520 95350
rect 205590 95150 205910 95350
rect 205980 95150 206020 95350
rect 206090 95150 206410 95350
rect 206480 95150 206520 95350
rect 206590 95150 206910 95350
rect 206980 95150 207020 95350
rect 207090 95150 207410 95350
rect 207480 95150 207520 95350
rect 207590 95150 207910 95350
rect 207980 95150 208000 95350
rect 196000 95140 208000 95150
rect 196140 95090 196360 95140
rect 196140 95020 196150 95090
rect 196350 95020 196360 95090
rect 196140 94980 196360 95020
rect 196140 94910 196150 94980
rect 196350 94910 196360 94980
rect 196140 94860 196360 94910
rect 196640 95090 196860 95140
rect 196640 95020 196650 95090
rect 196850 95020 196860 95090
rect 196640 94980 196860 95020
rect 196640 94910 196650 94980
rect 196850 94910 196860 94980
rect 196640 94860 196860 94910
rect 197140 95090 197360 95140
rect 197140 95020 197150 95090
rect 197350 95020 197360 95090
rect 197140 94980 197360 95020
rect 197140 94910 197150 94980
rect 197350 94910 197360 94980
rect 197140 94860 197360 94910
rect 197640 95090 197860 95140
rect 197640 95020 197650 95090
rect 197850 95020 197860 95090
rect 197640 94980 197860 95020
rect 197640 94910 197650 94980
rect 197850 94910 197860 94980
rect 197640 94860 197860 94910
rect 198140 95090 198360 95140
rect 198140 95020 198150 95090
rect 198350 95020 198360 95090
rect 198140 94980 198360 95020
rect 198140 94910 198150 94980
rect 198350 94910 198360 94980
rect 198140 94860 198360 94910
rect 198640 95090 198860 95140
rect 198640 95020 198650 95090
rect 198850 95020 198860 95090
rect 198640 94980 198860 95020
rect 198640 94910 198650 94980
rect 198850 94910 198860 94980
rect 198640 94860 198860 94910
rect 199140 95090 199360 95140
rect 199140 95020 199150 95090
rect 199350 95020 199360 95090
rect 199140 94980 199360 95020
rect 199140 94910 199150 94980
rect 199350 94910 199360 94980
rect 199140 94860 199360 94910
rect 199640 95090 199860 95140
rect 199640 95020 199650 95090
rect 199850 95020 199860 95090
rect 199640 94980 199860 95020
rect 199640 94910 199650 94980
rect 199850 94910 199860 94980
rect 199640 94860 199860 94910
rect 200140 95090 200360 95140
rect 200140 95020 200150 95090
rect 200350 95020 200360 95090
rect 200140 94980 200360 95020
rect 200140 94910 200150 94980
rect 200350 94910 200360 94980
rect 200140 94860 200360 94910
rect 200640 95090 200860 95140
rect 200640 95020 200650 95090
rect 200850 95020 200860 95090
rect 200640 94980 200860 95020
rect 200640 94910 200650 94980
rect 200850 94910 200860 94980
rect 200640 94860 200860 94910
rect 201140 95090 201360 95140
rect 201140 95020 201150 95090
rect 201350 95020 201360 95090
rect 201140 94980 201360 95020
rect 201140 94910 201150 94980
rect 201350 94910 201360 94980
rect 201140 94860 201360 94910
rect 201640 95090 201860 95140
rect 201640 95020 201650 95090
rect 201850 95020 201860 95090
rect 201640 94980 201860 95020
rect 201640 94910 201650 94980
rect 201850 94910 201860 94980
rect 201640 94860 201860 94910
rect 202140 95090 202360 95140
rect 202140 95020 202150 95090
rect 202350 95020 202360 95090
rect 202140 94980 202360 95020
rect 202140 94910 202150 94980
rect 202350 94910 202360 94980
rect 202140 94860 202360 94910
rect 202640 95090 202860 95140
rect 202640 95020 202650 95090
rect 202850 95020 202860 95090
rect 202640 94980 202860 95020
rect 202640 94910 202650 94980
rect 202850 94910 202860 94980
rect 202640 94860 202860 94910
rect 203140 95090 203360 95140
rect 203140 95020 203150 95090
rect 203350 95020 203360 95090
rect 203140 94980 203360 95020
rect 203140 94910 203150 94980
rect 203350 94910 203360 94980
rect 203140 94860 203360 94910
rect 203640 95090 203860 95140
rect 203640 95020 203650 95090
rect 203850 95020 203860 95090
rect 203640 94980 203860 95020
rect 203640 94910 203650 94980
rect 203850 94910 203860 94980
rect 203640 94860 203860 94910
rect 204140 95090 204360 95140
rect 204140 95020 204150 95090
rect 204350 95020 204360 95090
rect 204140 94980 204360 95020
rect 204140 94910 204150 94980
rect 204350 94910 204360 94980
rect 204140 94860 204360 94910
rect 204640 95090 204860 95140
rect 204640 95020 204650 95090
rect 204850 95020 204860 95090
rect 204640 94980 204860 95020
rect 204640 94910 204650 94980
rect 204850 94910 204860 94980
rect 204640 94860 204860 94910
rect 205140 95090 205360 95140
rect 205140 95020 205150 95090
rect 205350 95020 205360 95090
rect 205140 94980 205360 95020
rect 205140 94910 205150 94980
rect 205350 94910 205360 94980
rect 205140 94860 205360 94910
rect 205640 95090 205860 95140
rect 205640 95020 205650 95090
rect 205850 95020 205860 95090
rect 205640 94980 205860 95020
rect 205640 94910 205650 94980
rect 205850 94910 205860 94980
rect 205640 94860 205860 94910
rect 206140 95090 206360 95140
rect 206140 95020 206150 95090
rect 206350 95020 206360 95090
rect 206140 94980 206360 95020
rect 206140 94910 206150 94980
rect 206350 94910 206360 94980
rect 206140 94860 206360 94910
rect 206640 95090 206860 95140
rect 206640 95020 206650 95090
rect 206850 95020 206860 95090
rect 206640 94980 206860 95020
rect 206640 94910 206650 94980
rect 206850 94910 206860 94980
rect 206640 94860 206860 94910
rect 207140 95090 207360 95140
rect 207140 95020 207150 95090
rect 207350 95020 207360 95090
rect 207140 94980 207360 95020
rect 207140 94910 207150 94980
rect 207350 94910 207360 94980
rect 207140 94860 207360 94910
rect 207640 95090 207860 95140
rect 207640 95020 207650 95090
rect 207850 95020 207860 95090
rect 207640 94980 207860 95020
rect 207640 94910 207650 94980
rect 207850 94910 207860 94980
rect 207640 94860 207860 94910
rect 196000 94850 208000 94860
rect 196000 94650 196020 94850
rect 196090 94650 196410 94850
rect 196480 94650 196520 94850
rect 196590 94650 196910 94850
rect 196980 94650 197020 94850
rect 197090 94650 197410 94850
rect 197480 94650 197520 94850
rect 197590 94650 197910 94850
rect 197980 94650 198020 94850
rect 198090 94650 198410 94850
rect 198480 94650 198520 94850
rect 198590 94650 198910 94850
rect 198980 94650 199020 94850
rect 199090 94650 199410 94850
rect 199480 94650 199520 94850
rect 199590 94650 199910 94850
rect 199980 94650 200020 94850
rect 200090 94650 200410 94850
rect 200480 94650 200520 94850
rect 200590 94650 200910 94850
rect 200980 94650 201020 94850
rect 201090 94650 201410 94850
rect 201480 94650 201520 94850
rect 201590 94650 201910 94850
rect 201980 94650 202020 94850
rect 202090 94650 202410 94850
rect 202480 94650 202520 94850
rect 202590 94650 202910 94850
rect 202980 94650 203020 94850
rect 203090 94650 203410 94850
rect 203480 94650 203520 94850
rect 203590 94650 203910 94850
rect 203980 94650 204020 94850
rect 204090 94650 204410 94850
rect 204480 94650 204520 94850
rect 204590 94650 204910 94850
rect 204980 94650 205020 94850
rect 205090 94650 205410 94850
rect 205480 94650 205520 94850
rect 205590 94650 205910 94850
rect 205980 94650 206020 94850
rect 206090 94650 206410 94850
rect 206480 94650 206520 94850
rect 206590 94650 206910 94850
rect 206980 94650 207020 94850
rect 207090 94650 207410 94850
rect 207480 94650 207520 94850
rect 207590 94650 207910 94850
rect 207980 94650 208000 94850
rect 196000 94640 208000 94650
rect 196140 94590 196360 94640
rect 196140 94520 196150 94590
rect 196350 94520 196360 94590
rect 196140 94480 196360 94520
rect 196140 94410 196150 94480
rect 196350 94410 196360 94480
rect 196140 94360 196360 94410
rect 196640 94590 196860 94640
rect 196640 94520 196650 94590
rect 196850 94520 196860 94590
rect 196640 94480 196860 94520
rect 196640 94410 196650 94480
rect 196850 94410 196860 94480
rect 196640 94360 196860 94410
rect 197140 94590 197360 94640
rect 197140 94520 197150 94590
rect 197350 94520 197360 94590
rect 197140 94480 197360 94520
rect 197140 94410 197150 94480
rect 197350 94410 197360 94480
rect 197140 94360 197360 94410
rect 197640 94590 197860 94640
rect 197640 94520 197650 94590
rect 197850 94520 197860 94590
rect 197640 94480 197860 94520
rect 197640 94410 197650 94480
rect 197850 94410 197860 94480
rect 197640 94360 197860 94410
rect 198140 94590 198360 94640
rect 198140 94520 198150 94590
rect 198350 94520 198360 94590
rect 198140 94480 198360 94520
rect 198140 94410 198150 94480
rect 198350 94410 198360 94480
rect 198140 94360 198360 94410
rect 198640 94590 198860 94640
rect 198640 94520 198650 94590
rect 198850 94520 198860 94590
rect 198640 94480 198860 94520
rect 198640 94410 198650 94480
rect 198850 94410 198860 94480
rect 198640 94360 198860 94410
rect 199140 94590 199360 94640
rect 199140 94520 199150 94590
rect 199350 94520 199360 94590
rect 199140 94480 199360 94520
rect 199140 94410 199150 94480
rect 199350 94410 199360 94480
rect 199140 94360 199360 94410
rect 199640 94590 199860 94640
rect 199640 94520 199650 94590
rect 199850 94520 199860 94590
rect 199640 94480 199860 94520
rect 199640 94410 199650 94480
rect 199850 94410 199860 94480
rect 199640 94360 199860 94410
rect 200140 94590 200360 94640
rect 200140 94520 200150 94590
rect 200350 94520 200360 94590
rect 200140 94480 200360 94520
rect 200140 94410 200150 94480
rect 200350 94410 200360 94480
rect 200140 94360 200360 94410
rect 200640 94590 200860 94640
rect 200640 94520 200650 94590
rect 200850 94520 200860 94590
rect 200640 94480 200860 94520
rect 200640 94410 200650 94480
rect 200850 94410 200860 94480
rect 200640 94360 200860 94410
rect 201140 94590 201360 94640
rect 201140 94520 201150 94590
rect 201350 94520 201360 94590
rect 201140 94480 201360 94520
rect 201140 94410 201150 94480
rect 201350 94410 201360 94480
rect 201140 94360 201360 94410
rect 201640 94590 201860 94640
rect 201640 94520 201650 94590
rect 201850 94520 201860 94590
rect 201640 94480 201860 94520
rect 201640 94410 201650 94480
rect 201850 94410 201860 94480
rect 201640 94360 201860 94410
rect 202140 94590 202360 94640
rect 202140 94520 202150 94590
rect 202350 94520 202360 94590
rect 202140 94480 202360 94520
rect 202140 94410 202150 94480
rect 202350 94410 202360 94480
rect 202140 94360 202360 94410
rect 202640 94590 202860 94640
rect 202640 94520 202650 94590
rect 202850 94520 202860 94590
rect 202640 94480 202860 94520
rect 202640 94410 202650 94480
rect 202850 94410 202860 94480
rect 202640 94360 202860 94410
rect 203140 94590 203360 94640
rect 203140 94520 203150 94590
rect 203350 94520 203360 94590
rect 203140 94480 203360 94520
rect 203140 94410 203150 94480
rect 203350 94410 203360 94480
rect 203140 94360 203360 94410
rect 203640 94590 203860 94640
rect 203640 94520 203650 94590
rect 203850 94520 203860 94590
rect 203640 94480 203860 94520
rect 203640 94410 203650 94480
rect 203850 94410 203860 94480
rect 203640 94360 203860 94410
rect 204140 94590 204360 94640
rect 204140 94520 204150 94590
rect 204350 94520 204360 94590
rect 204140 94480 204360 94520
rect 204140 94410 204150 94480
rect 204350 94410 204360 94480
rect 204140 94360 204360 94410
rect 204640 94590 204860 94640
rect 204640 94520 204650 94590
rect 204850 94520 204860 94590
rect 204640 94480 204860 94520
rect 204640 94410 204650 94480
rect 204850 94410 204860 94480
rect 204640 94360 204860 94410
rect 205140 94590 205360 94640
rect 205140 94520 205150 94590
rect 205350 94520 205360 94590
rect 205140 94480 205360 94520
rect 205140 94410 205150 94480
rect 205350 94410 205360 94480
rect 205140 94360 205360 94410
rect 205640 94590 205860 94640
rect 205640 94520 205650 94590
rect 205850 94520 205860 94590
rect 205640 94480 205860 94520
rect 205640 94410 205650 94480
rect 205850 94410 205860 94480
rect 205640 94360 205860 94410
rect 206140 94590 206360 94640
rect 206140 94520 206150 94590
rect 206350 94520 206360 94590
rect 206140 94480 206360 94520
rect 206140 94410 206150 94480
rect 206350 94410 206360 94480
rect 206140 94360 206360 94410
rect 206640 94590 206860 94640
rect 206640 94520 206650 94590
rect 206850 94520 206860 94590
rect 206640 94480 206860 94520
rect 206640 94410 206650 94480
rect 206850 94410 206860 94480
rect 206640 94360 206860 94410
rect 207140 94590 207360 94640
rect 207140 94520 207150 94590
rect 207350 94520 207360 94590
rect 207140 94480 207360 94520
rect 207140 94410 207150 94480
rect 207350 94410 207360 94480
rect 207140 94360 207360 94410
rect 207640 94590 207860 94640
rect 207640 94520 207650 94590
rect 207850 94520 207860 94590
rect 207640 94480 207860 94520
rect 207640 94410 207650 94480
rect 207850 94410 207860 94480
rect 207640 94360 207860 94410
rect 196000 94350 208000 94360
rect 196000 94150 196020 94350
rect 196090 94150 196410 94350
rect 196480 94150 196520 94350
rect 196590 94150 196910 94350
rect 196980 94150 197020 94350
rect 197090 94150 197410 94350
rect 197480 94150 197520 94350
rect 197590 94150 197910 94350
rect 197980 94150 198020 94350
rect 198090 94150 198410 94350
rect 198480 94150 198520 94350
rect 198590 94150 198910 94350
rect 198980 94150 199020 94350
rect 199090 94150 199410 94350
rect 199480 94150 199520 94350
rect 199590 94150 199910 94350
rect 199980 94150 200020 94350
rect 200090 94150 200410 94350
rect 200480 94150 200520 94350
rect 200590 94150 200910 94350
rect 200980 94150 201020 94350
rect 201090 94150 201410 94350
rect 201480 94150 201520 94350
rect 201590 94150 201910 94350
rect 201980 94150 202020 94350
rect 202090 94150 202410 94350
rect 202480 94150 202520 94350
rect 202590 94150 202910 94350
rect 202980 94150 203020 94350
rect 203090 94150 203410 94350
rect 203480 94150 203520 94350
rect 203590 94150 203910 94350
rect 203980 94150 204020 94350
rect 204090 94150 204410 94350
rect 204480 94150 204520 94350
rect 204590 94150 204910 94350
rect 204980 94150 205020 94350
rect 205090 94150 205410 94350
rect 205480 94150 205520 94350
rect 205590 94150 205910 94350
rect 205980 94150 206020 94350
rect 206090 94150 206410 94350
rect 206480 94150 206520 94350
rect 206590 94150 206910 94350
rect 206980 94150 207020 94350
rect 207090 94150 207410 94350
rect 207480 94150 207520 94350
rect 207590 94150 207910 94350
rect 207980 94150 208000 94350
rect 196000 94140 208000 94150
rect 196140 94090 196360 94140
rect 196140 94020 196150 94090
rect 196350 94020 196360 94090
rect 196140 93980 196360 94020
rect 196140 93910 196150 93980
rect 196350 93910 196360 93980
rect 196140 93860 196360 93910
rect 196640 94090 196860 94140
rect 196640 94020 196650 94090
rect 196850 94020 196860 94090
rect 196640 93980 196860 94020
rect 196640 93910 196650 93980
rect 196850 93910 196860 93980
rect 196640 93860 196860 93910
rect 197140 94090 197360 94140
rect 197140 94020 197150 94090
rect 197350 94020 197360 94090
rect 197140 93980 197360 94020
rect 197140 93910 197150 93980
rect 197350 93910 197360 93980
rect 197140 93860 197360 93910
rect 197640 94090 197860 94140
rect 197640 94020 197650 94090
rect 197850 94020 197860 94090
rect 197640 93980 197860 94020
rect 197640 93910 197650 93980
rect 197850 93910 197860 93980
rect 197640 93860 197860 93910
rect 198140 94090 198360 94140
rect 198140 94020 198150 94090
rect 198350 94020 198360 94090
rect 198140 93980 198360 94020
rect 198140 93910 198150 93980
rect 198350 93910 198360 93980
rect 198140 93860 198360 93910
rect 198640 94090 198860 94140
rect 198640 94020 198650 94090
rect 198850 94020 198860 94090
rect 198640 93980 198860 94020
rect 198640 93910 198650 93980
rect 198850 93910 198860 93980
rect 198640 93860 198860 93910
rect 199140 94090 199360 94140
rect 199140 94020 199150 94090
rect 199350 94020 199360 94090
rect 199140 93980 199360 94020
rect 199140 93910 199150 93980
rect 199350 93910 199360 93980
rect 199140 93860 199360 93910
rect 199640 94090 199860 94140
rect 199640 94020 199650 94090
rect 199850 94020 199860 94090
rect 199640 93980 199860 94020
rect 199640 93910 199650 93980
rect 199850 93910 199860 93980
rect 199640 93860 199860 93910
rect 200140 94090 200360 94140
rect 200140 94020 200150 94090
rect 200350 94020 200360 94090
rect 200140 93980 200360 94020
rect 200140 93910 200150 93980
rect 200350 93910 200360 93980
rect 200140 93860 200360 93910
rect 200640 94090 200860 94140
rect 200640 94020 200650 94090
rect 200850 94020 200860 94090
rect 200640 93980 200860 94020
rect 200640 93910 200650 93980
rect 200850 93910 200860 93980
rect 200640 93860 200860 93910
rect 201140 94090 201360 94140
rect 201140 94020 201150 94090
rect 201350 94020 201360 94090
rect 201140 93980 201360 94020
rect 201140 93910 201150 93980
rect 201350 93910 201360 93980
rect 201140 93860 201360 93910
rect 201640 94090 201860 94140
rect 201640 94020 201650 94090
rect 201850 94020 201860 94090
rect 201640 93980 201860 94020
rect 201640 93910 201650 93980
rect 201850 93910 201860 93980
rect 201640 93860 201860 93910
rect 202140 94090 202360 94140
rect 202140 94020 202150 94090
rect 202350 94020 202360 94090
rect 202140 93980 202360 94020
rect 202140 93910 202150 93980
rect 202350 93910 202360 93980
rect 202140 93860 202360 93910
rect 202640 94090 202860 94140
rect 202640 94020 202650 94090
rect 202850 94020 202860 94090
rect 202640 93980 202860 94020
rect 202640 93910 202650 93980
rect 202850 93910 202860 93980
rect 202640 93860 202860 93910
rect 203140 94090 203360 94140
rect 203140 94020 203150 94090
rect 203350 94020 203360 94090
rect 203140 93980 203360 94020
rect 203140 93910 203150 93980
rect 203350 93910 203360 93980
rect 203140 93860 203360 93910
rect 203640 94090 203860 94140
rect 203640 94020 203650 94090
rect 203850 94020 203860 94090
rect 203640 93980 203860 94020
rect 203640 93910 203650 93980
rect 203850 93910 203860 93980
rect 203640 93860 203860 93910
rect 204140 94090 204360 94140
rect 204140 94020 204150 94090
rect 204350 94020 204360 94090
rect 204140 93980 204360 94020
rect 204140 93910 204150 93980
rect 204350 93910 204360 93980
rect 204140 93860 204360 93910
rect 204640 94090 204860 94140
rect 204640 94020 204650 94090
rect 204850 94020 204860 94090
rect 204640 93980 204860 94020
rect 204640 93910 204650 93980
rect 204850 93910 204860 93980
rect 204640 93860 204860 93910
rect 205140 94090 205360 94140
rect 205140 94020 205150 94090
rect 205350 94020 205360 94090
rect 205140 93980 205360 94020
rect 205140 93910 205150 93980
rect 205350 93910 205360 93980
rect 205140 93860 205360 93910
rect 205640 94090 205860 94140
rect 205640 94020 205650 94090
rect 205850 94020 205860 94090
rect 205640 93980 205860 94020
rect 205640 93910 205650 93980
rect 205850 93910 205860 93980
rect 205640 93860 205860 93910
rect 206140 94090 206360 94140
rect 206140 94020 206150 94090
rect 206350 94020 206360 94090
rect 206140 93980 206360 94020
rect 206140 93910 206150 93980
rect 206350 93910 206360 93980
rect 206140 93860 206360 93910
rect 206640 94090 206860 94140
rect 206640 94020 206650 94090
rect 206850 94020 206860 94090
rect 206640 93980 206860 94020
rect 206640 93910 206650 93980
rect 206850 93910 206860 93980
rect 206640 93860 206860 93910
rect 207140 94090 207360 94140
rect 207140 94020 207150 94090
rect 207350 94020 207360 94090
rect 207140 93980 207360 94020
rect 207140 93910 207150 93980
rect 207350 93910 207360 93980
rect 207140 93860 207360 93910
rect 207640 94090 207860 94140
rect 207640 94020 207650 94090
rect 207850 94020 207860 94090
rect 207640 93980 207860 94020
rect 207640 93910 207650 93980
rect 207850 93910 207860 93980
rect 207640 93860 207860 93910
rect 196000 93850 208000 93860
rect 196000 93650 196020 93850
rect 196090 93650 196410 93850
rect 196480 93650 196520 93850
rect 196590 93650 196910 93850
rect 196980 93650 197020 93850
rect 197090 93650 197410 93850
rect 197480 93650 197520 93850
rect 197590 93650 197910 93850
rect 197980 93650 198020 93850
rect 198090 93650 198410 93850
rect 198480 93650 198520 93850
rect 198590 93650 198910 93850
rect 198980 93650 199020 93850
rect 199090 93650 199410 93850
rect 199480 93650 199520 93850
rect 199590 93650 199910 93850
rect 199980 93650 200020 93850
rect 200090 93650 200410 93850
rect 200480 93650 200520 93850
rect 200590 93650 200910 93850
rect 200980 93650 201020 93850
rect 201090 93650 201410 93850
rect 201480 93650 201520 93850
rect 201590 93650 201910 93850
rect 201980 93650 202020 93850
rect 202090 93650 202410 93850
rect 202480 93650 202520 93850
rect 202590 93650 202910 93850
rect 202980 93650 203020 93850
rect 203090 93650 203410 93850
rect 203480 93650 203520 93850
rect 203590 93650 203910 93850
rect 203980 93650 204020 93850
rect 204090 93650 204410 93850
rect 204480 93650 204520 93850
rect 204590 93650 204910 93850
rect 204980 93650 205020 93850
rect 205090 93650 205410 93850
rect 205480 93650 205520 93850
rect 205590 93650 205910 93850
rect 205980 93650 206020 93850
rect 206090 93650 206410 93850
rect 206480 93650 206520 93850
rect 206590 93650 206910 93850
rect 206980 93650 207020 93850
rect 207090 93650 207410 93850
rect 207480 93650 207520 93850
rect 207590 93650 207910 93850
rect 207980 93650 208000 93850
rect 196000 93640 208000 93650
rect 196140 93590 196360 93640
rect 196140 93520 196150 93590
rect 196350 93520 196360 93590
rect 196140 93480 196360 93520
rect 196140 93410 196150 93480
rect 196350 93410 196360 93480
rect 196140 93360 196360 93410
rect 196640 93590 196860 93640
rect 196640 93520 196650 93590
rect 196850 93520 196860 93590
rect 196640 93480 196860 93520
rect 196640 93410 196650 93480
rect 196850 93410 196860 93480
rect 196640 93360 196860 93410
rect 197140 93590 197360 93640
rect 197140 93520 197150 93590
rect 197350 93520 197360 93590
rect 197140 93480 197360 93520
rect 197140 93410 197150 93480
rect 197350 93410 197360 93480
rect 197140 93360 197360 93410
rect 197640 93590 197860 93640
rect 197640 93520 197650 93590
rect 197850 93520 197860 93590
rect 197640 93480 197860 93520
rect 197640 93410 197650 93480
rect 197850 93410 197860 93480
rect 197640 93360 197860 93410
rect 198140 93590 198360 93640
rect 198140 93520 198150 93590
rect 198350 93520 198360 93590
rect 198140 93480 198360 93520
rect 198140 93410 198150 93480
rect 198350 93410 198360 93480
rect 198140 93360 198360 93410
rect 198640 93590 198860 93640
rect 198640 93520 198650 93590
rect 198850 93520 198860 93590
rect 198640 93480 198860 93520
rect 198640 93410 198650 93480
rect 198850 93410 198860 93480
rect 198640 93360 198860 93410
rect 199140 93590 199360 93640
rect 199140 93520 199150 93590
rect 199350 93520 199360 93590
rect 199140 93480 199360 93520
rect 199140 93410 199150 93480
rect 199350 93410 199360 93480
rect 199140 93360 199360 93410
rect 199640 93590 199860 93640
rect 199640 93520 199650 93590
rect 199850 93520 199860 93590
rect 199640 93480 199860 93520
rect 199640 93410 199650 93480
rect 199850 93410 199860 93480
rect 199640 93360 199860 93410
rect 200140 93590 200360 93640
rect 200140 93520 200150 93590
rect 200350 93520 200360 93590
rect 200140 93480 200360 93520
rect 200140 93410 200150 93480
rect 200350 93410 200360 93480
rect 200140 93360 200360 93410
rect 200640 93590 200860 93640
rect 200640 93520 200650 93590
rect 200850 93520 200860 93590
rect 200640 93480 200860 93520
rect 200640 93410 200650 93480
rect 200850 93410 200860 93480
rect 200640 93360 200860 93410
rect 201140 93590 201360 93640
rect 201140 93520 201150 93590
rect 201350 93520 201360 93590
rect 201140 93480 201360 93520
rect 201140 93410 201150 93480
rect 201350 93410 201360 93480
rect 201140 93360 201360 93410
rect 201640 93590 201860 93640
rect 201640 93520 201650 93590
rect 201850 93520 201860 93590
rect 201640 93480 201860 93520
rect 201640 93410 201650 93480
rect 201850 93410 201860 93480
rect 201640 93360 201860 93410
rect 202140 93590 202360 93640
rect 202140 93520 202150 93590
rect 202350 93520 202360 93590
rect 202140 93480 202360 93520
rect 202140 93410 202150 93480
rect 202350 93410 202360 93480
rect 202140 93360 202360 93410
rect 202640 93590 202860 93640
rect 202640 93520 202650 93590
rect 202850 93520 202860 93590
rect 202640 93480 202860 93520
rect 202640 93410 202650 93480
rect 202850 93410 202860 93480
rect 202640 93360 202860 93410
rect 203140 93590 203360 93640
rect 203140 93520 203150 93590
rect 203350 93520 203360 93590
rect 203140 93480 203360 93520
rect 203140 93410 203150 93480
rect 203350 93410 203360 93480
rect 203140 93360 203360 93410
rect 203640 93590 203860 93640
rect 203640 93520 203650 93590
rect 203850 93520 203860 93590
rect 203640 93480 203860 93520
rect 203640 93410 203650 93480
rect 203850 93410 203860 93480
rect 203640 93360 203860 93410
rect 204140 93590 204360 93640
rect 204140 93520 204150 93590
rect 204350 93520 204360 93590
rect 204140 93480 204360 93520
rect 204140 93410 204150 93480
rect 204350 93410 204360 93480
rect 204140 93360 204360 93410
rect 204640 93590 204860 93640
rect 204640 93520 204650 93590
rect 204850 93520 204860 93590
rect 204640 93480 204860 93520
rect 204640 93410 204650 93480
rect 204850 93410 204860 93480
rect 204640 93360 204860 93410
rect 205140 93590 205360 93640
rect 205140 93520 205150 93590
rect 205350 93520 205360 93590
rect 205140 93480 205360 93520
rect 205140 93410 205150 93480
rect 205350 93410 205360 93480
rect 205140 93360 205360 93410
rect 205640 93590 205860 93640
rect 205640 93520 205650 93590
rect 205850 93520 205860 93590
rect 205640 93480 205860 93520
rect 205640 93410 205650 93480
rect 205850 93410 205860 93480
rect 205640 93360 205860 93410
rect 206140 93590 206360 93640
rect 206140 93520 206150 93590
rect 206350 93520 206360 93590
rect 206140 93480 206360 93520
rect 206140 93410 206150 93480
rect 206350 93410 206360 93480
rect 206140 93360 206360 93410
rect 206640 93590 206860 93640
rect 206640 93520 206650 93590
rect 206850 93520 206860 93590
rect 206640 93480 206860 93520
rect 206640 93410 206650 93480
rect 206850 93410 206860 93480
rect 206640 93360 206860 93410
rect 207140 93590 207360 93640
rect 207140 93520 207150 93590
rect 207350 93520 207360 93590
rect 207140 93480 207360 93520
rect 207140 93410 207150 93480
rect 207350 93410 207360 93480
rect 207140 93360 207360 93410
rect 207640 93590 207860 93640
rect 207640 93520 207650 93590
rect 207850 93520 207860 93590
rect 207640 93480 207860 93520
rect 207640 93410 207650 93480
rect 207850 93410 207860 93480
rect 207640 93360 207860 93410
rect 196000 93350 208000 93360
rect 196000 93150 196020 93350
rect 196090 93150 196410 93350
rect 196480 93150 196520 93350
rect 196590 93150 196910 93350
rect 196980 93150 197020 93350
rect 197090 93150 197410 93350
rect 197480 93150 197520 93350
rect 197590 93150 197910 93350
rect 197980 93150 198020 93350
rect 198090 93150 198410 93350
rect 198480 93150 198520 93350
rect 198590 93150 198910 93350
rect 198980 93150 199020 93350
rect 199090 93150 199410 93350
rect 199480 93150 199520 93350
rect 199590 93150 199910 93350
rect 199980 93150 200020 93350
rect 200090 93150 200410 93350
rect 200480 93150 200520 93350
rect 200590 93150 200910 93350
rect 200980 93150 201020 93350
rect 201090 93150 201410 93350
rect 201480 93150 201520 93350
rect 201590 93150 201910 93350
rect 201980 93150 202020 93350
rect 202090 93150 202410 93350
rect 202480 93150 202520 93350
rect 202590 93150 202910 93350
rect 202980 93150 203020 93350
rect 203090 93150 203410 93350
rect 203480 93150 203520 93350
rect 203590 93150 203910 93350
rect 203980 93150 204020 93350
rect 204090 93150 204410 93350
rect 204480 93150 204520 93350
rect 204590 93150 204910 93350
rect 204980 93150 205020 93350
rect 205090 93150 205410 93350
rect 205480 93150 205520 93350
rect 205590 93150 205910 93350
rect 205980 93150 206020 93350
rect 206090 93150 206410 93350
rect 206480 93150 206520 93350
rect 206590 93150 206910 93350
rect 206980 93150 207020 93350
rect 207090 93150 207410 93350
rect 207480 93150 207520 93350
rect 207590 93150 207910 93350
rect 207980 93150 208000 93350
rect 196000 93140 208000 93150
rect 196140 93090 196360 93140
rect 196140 93020 196150 93090
rect 196350 93020 196360 93090
rect 196140 92980 196360 93020
rect 196140 92910 196150 92980
rect 196350 92910 196360 92980
rect 196140 92860 196360 92910
rect 196640 93090 196860 93140
rect 196640 93020 196650 93090
rect 196850 93020 196860 93090
rect 196640 92980 196860 93020
rect 196640 92910 196650 92980
rect 196850 92910 196860 92980
rect 196640 92860 196860 92910
rect 197140 93090 197360 93140
rect 197140 93020 197150 93090
rect 197350 93020 197360 93090
rect 197140 92980 197360 93020
rect 197140 92910 197150 92980
rect 197350 92910 197360 92980
rect 197140 92860 197360 92910
rect 197640 93090 197860 93140
rect 197640 93020 197650 93090
rect 197850 93020 197860 93090
rect 197640 92980 197860 93020
rect 197640 92910 197650 92980
rect 197850 92910 197860 92980
rect 197640 92860 197860 92910
rect 198140 93090 198360 93140
rect 198140 93020 198150 93090
rect 198350 93020 198360 93090
rect 198140 92980 198360 93020
rect 198140 92910 198150 92980
rect 198350 92910 198360 92980
rect 198140 92860 198360 92910
rect 198640 93090 198860 93140
rect 198640 93020 198650 93090
rect 198850 93020 198860 93090
rect 198640 92980 198860 93020
rect 198640 92910 198650 92980
rect 198850 92910 198860 92980
rect 198640 92860 198860 92910
rect 199140 93090 199360 93140
rect 199140 93020 199150 93090
rect 199350 93020 199360 93090
rect 199140 92980 199360 93020
rect 199140 92910 199150 92980
rect 199350 92910 199360 92980
rect 199140 92860 199360 92910
rect 199640 93090 199860 93140
rect 199640 93020 199650 93090
rect 199850 93020 199860 93090
rect 199640 92980 199860 93020
rect 199640 92910 199650 92980
rect 199850 92910 199860 92980
rect 199640 92860 199860 92910
rect 200140 93090 200360 93140
rect 200140 93020 200150 93090
rect 200350 93020 200360 93090
rect 200140 92980 200360 93020
rect 200140 92910 200150 92980
rect 200350 92910 200360 92980
rect 200140 92860 200360 92910
rect 200640 93090 200860 93140
rect 200640 93020 200650 93090
rect 200850 93020 200860 93090
rect 200640 92980 200860 93020
rect 200640 92910 200650 92980
rect 200850 92910 200860 92980
rect 200640 92860 200860 92910
rect 201140 93090 201360 93140
rect 201140 93020 201150 93090
rect 201350 93020 201360 93090
rect 201140 92980 201360 93020
rect 201140 92910 201150 92980
rect 201350 92910 201360 92980
rect 201140 92860 201360 92910
rect 201640 93090 201860 93140
rect 201640 93020 201650 93090
rect 201850 93020 201860 93090
rect 201640 92980 201860 93020
rect 201640 92910 201650 92980
rect 201850 92910 201860 92980
rect 201640 92860 201860 92910
rect 202140 93090 202360 93140
rect 202140 93020 202150 93090
rect 202350 93020 202360 93090
rect 202140 92980 202360 93020
rect 202140 92910 202150 92980
rect 202350 92910 202360 92980
rect 202140 92860 202360 92910
rect 202640 93090 202860 93140
rect 202640 93020 202650 93090
rect 202850 93020 202860 93090
rect 202640 92980 202860 93020
rect 202640 92910 202650 92980
rect 202850 92910 202860 92980
rect 202640 92860 202860 92910
rect 203140 93090 203360 93140
rect 203140 93020 203150 93090
rect 203350 93020 203360 93090
rect 203140 92980 203360 93020
rect 203140 92910 203150 92980
rect 203350 92910 203360 92980
rect 203140 92860 203360 92910
rect 203640 93090 203860 93140
rect 203640 93020 203650 93090
rect 203850 93020 203860 93090
rect 203640 92980 203860 93020
rect 203640 92910 203650 92980
rect 203850 92910 203860 92980
rect 203640 92860 203860 92910
rect 204140 93090 204360 93140
rect 204140 93020 204150 93090
rect 204350 93020 204360 93090
rect 204140 92980 204360 93020
rect 204140 92910 204150 92980
rect 204350 92910 204360 92980
rect 204140 92860 204360 92910
rect 204640 93090 204860 93140
rect 204640 93020 204650 93090
rect 204850 93020 204860 93090
rect 204640 92980 204860 93020
rect 204640 92910 204650 92980
rect 204850 92910 204860 92980
rect 204640 92860 204860 92910
rect 205140 93090 205360 93140
rect 205140 93020 205150 93090
rect 205350 93020 205360 93090
rect 205140 92980 205360 93020
rect 205140 92910 205150 92980
rect 205350 92910 205360 92980
rect 205140 92860 205360 92910
rect 205640 93090 205860 93140
rect 205640 93020 205650 93090
rect 205850 93020 205860 93090
rect 205640 92980 205860 93020
rect 205640 92910 205650 92980
rect 205850 92910 205860 92980
rect 205640 92860 205860 92910
rect 206140 93090 206360 93140
rect 206140 93020 206150 93090
rect 206350 93020 206360 93090
rect 206140 92980 206360 93020
rect 206140 92910 206150 92980
rect 206350 92910 206360 92980
rect 206140 92860 206360 92910
rect 206640 93090 206860 93140
rect 206640 93020 206650 93090
rect 206850 93020 206860 93090
rect 206640 92980 206860 93020
rect 206640 92910 206650 92980
rect 206850 92910 206860 92980
rect 206640 92860 206860 92910
rect 207140 93090 207360 93140
rect 207140 93020 207150 93090
rect 207350 93020 207360 93090
rect 207140 92980 207360 93020
rect 207140 92910 207150 92980
rect 207350 92910 207360 92980
rect 207140 92860 207360 92910
rect 207640 93090 207860 93140
rect 207640 93020 207650 93090
rect 207850 93020 207860 93090
rect 207640 92980 207860 93020
rect 207640 92910 207650 92980
rect 207850 92910 207860 92980
rect 207640 92860 207860 92910
rect 196000 92850 208000 92860
rect 196000 92650 196020 92850
rect 196090 92650 196410 92850
rect 196480 92650 196520 92850
rect 196590 92650 196910 92850
rect 196980 92650 197020 92850
rect 197090 92650 197410 92850
rect 197480 92650 197520 92850
rect 197590 92650 197910 92850
rect 197980 92650 198020 92850
rect 198090 92650 198410 92850
rect 198480 92650 198520 92850
rect 198590 92650 198910 92850
rect 198980 92650 199020 92850
rect 199090 92650 199410 92850
rect 199480 92650 199520 92850
rect 199590 92650 199910 92850
rect 199980 92650 200020 92850
rect 200090 92650 200410 92850
rect 200480 92650 200520 92850
rect 200590 92650 200910 92850
rect 200980 92650 201020 92850
rect 201090 92650 201410 92850
rect 201480 92650 201520 92850
rect 201590 92650 201910 92850
rect 201980 92650 202020 92850
rect 202090 92650 202410 92850
rect 202480 92650 202520 92850
rect 202590 92650 202910 92850
rect 202980 92650 203020 92850
rect 203090 92650 203410 92850
rect 203480 92650 203520 92850
rect 203590 92650 203910 92850
rect 203980 92650 204020 92850
rect 204090 92650 204410 92850
rect 204480 92650 204520 92850
rect 204590 92650 204910 92850
rect 204980 92650 205020 92850
rect 205090 92650 205410 92850
rect 205480 92650 205520 92850
rect 205590 92650 205910 92850
rect 205980 92650 206020 92850
rect 206090 92650 206410 92850
rect 206480 92650 206520 92850
rect 206590 92650 206910 92850
rect 206980 92650 207020 92850
rect 207090 92650 207410 92850
rect 207480 92650 207520 92850
rect 207590 92650 207910 92850
rect 207980 92650 208000 92850
rect 196000 92640 208000 92650
rect 196140 92590 196360 92640
rect 196140 92520 196150 92590
rect 196350 92520 196360 92590
rect 196140 92480 196360 92520
rect 196140 92410 196150 92480
rect 196350 92410 196360 92480
rect 196140 92360 196360 92410
rect 196640 92590 196860 92640
rect 196640 92520 196650 92590
rect 196850 92520 196860 92590
rect 196640 92480 196860 92520
rect 196640 92410 196650 92480
rect 196850 92410 196860 92480
rect 196640 92360 196860 92410
rect 197140 92590 197360 92640
rect 197140 92520 197150 92590
rect 197350 92520 197360 92590
rect 197140 92480 197360 92520
rect 197140 92410 197150 92480
rect 197350 92410 197360 92480
rect 197140 92360 197360 92410
rect 197640 92590 197860 92640
rect 197640 92520 197650 92590
rect 197850 92520 197860 92590
rect 197640 92480 197860 92520
rect 197640 92410 197650 92480
rect 197850 92410 197860 92480
rect 197640 92360 197860 92410
rect 198140 92590 198360 92640
rect 198140 92520 198150 92590
rect 198350 92520 198360 92590
rect 198140 92480 198360 92520
rect 198140 92410 198150 92480
rect 198350 92410 198360 92480
rect 198140 92360 198360 92410
rect 198640 92590 198860 92640
rect 198640 92520 198650 92590
rect 198850 92520 198860 92590
rect 198640 92480 198860 92520
rect 198640 92410 198650 92480
rect 198850 92410 198860 92480
rect 198640 92360 198860 92410
rect 199140 92590 199360 92640
rect 199140 92520 199150 92590
rect 199350 92520 199360 92590
rect 199140 92480 199360 92520
rect 199140 92410 199150 92480
rect 199350 92410 199360 92480
rect 199140 92360 199360 92410
rect 199640 92590 199860 92640
rect 199640 92520 199650 92590
rect 199850 92520 199860 92590
rect 199640 92480 199860 92520
rect 199640 92410 199650 92480
rect 199850 92410 199860 92480
rect 199640 92360 199860 92410
rect 200140 92590 200360 92640
rect 200140 92520 200150 92590
rect 200350 92520 200360 92590
rect 200140 92480 200360 92520
rect 200140 92410 200150 92480
rect 200350 92410 200360 92480
rect 200140 92360 200360 92410
rect 200640 92590 200860 92640
rect 200640 92520 200650 92590
rect 200850 92520 200860 92590
rect 200640 92480 200860 92520
rect 200640 92410 200650 92480
rect 200850 92410 200860 92480
rect 200640 92360 200860 92410
rect 201140 92590 201360 92640
rect 201140 92520 201150 92590
rect 201350 92520 201360 92590
rect 201140 92480 201360 92520
rect 201140 92410 201150 92480
rect 201350 92410 201360 92480
rect 201140 92360 201360 92410
rect 201640 92590 201860 92640
rect 201640 92520 201650 92590
rect 201850 92520 201860 92590
rect 201640 92480 201860 92520
rect 201640 92410 201650 92480
rect 201850 92410 201860 92480
rect 201640 92360 201860 92410
rect 202140 92590 202360 92640
rect 202140 92520 202150 92590
rect 202350 92520 202360 92590
rect 202140 92480 202360 92520
rect 202140 92410 202150 92480
rect 202350 92410 202360 92480
rect 202140 92360 202360 92410
rect 202640 92590 202860 92640
rect 202640 92520 202650 92590
rect 202850 92520 202860 92590
rect 202640 92480 202860 92520
rect 202640 92410 202650 92480
rect 202850 92410 202860 92480
rect 202640 92360 202860 92410
rect 203140 92590 203360 92640
rect 203140 92520 203150 92590
rect 203350 92520 203360 92590
rect 203140 92480 203360 92520
rect 203140 92410 203150 92480
rect 203350 92410 203360 92480
rect 203140 92360 203360 92410
rect 203640 92590 203860 92640
rect 203640 92520 203650 92590
rect 203850 92520 203860 92590
rect 203640 92480 203860 92520
rect 203640 92410 203650 92480
rect 203850 92410 203860 92480
rect 203640 92360 203860 92410
rect 204140 92590 204360 92640
rect 204140 92520 204150 92590
rect 204350 92520 204360 92590
rect 204140 92480 204360 92520
rect 204140 92410 204150 92480
rect 204350 92410 204360 92480
rect 204140 92360 204360 92410
rect 204640 92590 204860 92640
rect 204640 92520 204650 92590
rect 204850 92520 204860 92590
rect 204640 92480 204860 92520
rect 204640 92410 204650 92480
rect 204850 92410 204860 92480
rect 204640 92360 204860 92410
rect 205140 92590 205360 92640
rect 205140 92520 205150 92590
rect 205350 92520 205360 92590
rect 205140 92480 205360 92520
rect 205140 92410 205150 92480
rect 205350 92410 205360 92480
rect 205140 92360 205360 92410
rect 205640 92590 205860 92640
rect 205640 92520 205650 92590
rect 205850 92520 205860 92590
rect 205640 92480 205860 92520
rect 205640 92410 205650 92480
rect 205850 92410 205860 92480
rect 205640 92360 205860 92410
rect 206140 92590 206360 92640
rect 206140 92520 206150 92590
rect 206350 92520 206360 92590
rect 206140 92480 206360 92520
rect 206140 92410 206150 92480
rect 206350 92410 206360 92480
rect 206140 92360 206360 92410
rect 206640 92590 206860 92640
rect 206640 92520 206650 92590
rect 206850 92520 206860 92590
rect 206640 92480 206860 92520
rect 206640 92410 206650 92480
rect 206850 92410 206860 92480
rect 206640 92360 206860 92410
rect 207140 92590 207360 92640
rect 207140 92520 207150 92590
rect 207350 92520 207360 92590
rect 207140 92480 207360 92520
rect 207140 92410 207150 92480
rect 207350 92410 207360 92480
rect 207140 92360 207360 92410
rect 207640 92590 207860 92640
rect 207640 92520 207650 92590
rect 207850 92520 207860 92590
rect 207640 92480 207860 92520
rect 207640 92410 207650 92480
rect 207850 92410 207860 92480
rect 207640 92360 207860 92410
rect 196000 92350 208000 92360
rect 196000 92150 196020 92350
rect 196090 92150 196410 92350
rect 196480 92150 196520 92350
rect 196590 92150 196910 92350
rect 196980 92150 197020 92350
rect 197090 92150 197410 92350
rect 197480 92150 197520 92350
rect 197590 92150 197910 92350
rect 197980 92150 198020 92350
rect 198090 92150 198410 92350
rect 198480 92150 198520 92350
rect 198590 92150 198910 92350
rect 198980 92150 199020 92350
rect 199090 92150 199410 92350
rect 199480 92150 199520 92350
rect 199590 92150 199910 92350
rect 199980 92150 200020 92350
rect 200090 92150 200410 92350
rect 200480 92150 200520 92350
rect 200590 92150 200910 92350
rect 200980 92150 201020 92350
rect 201090 92150 201410 92350
rect 201480 92150 201520 92350
rect 201590 92150 201910 92350
rect 201980 92150 202020 92350
rect 202090 92150 202410 92350
rect 202480 92150 202520 92350
rect 202590 92150 202910 92350
rect 202980 92150 203020 92350
rect 203090 92150 203410 92350
rect 203480 92150 203520 92350
rect 203590 92150 203910 92350
rect 203980 92150 204020 92350
rect 204090 92150 204410 92350
rect 204480 92150 204520 92350
rect 204590 92150 204910 92350
rect 204980 92150 205020 92350
rect 205090 92150 205410 92350
rect 205480 92150 205520 92350
rect 205590 92150 205910 92350
rect 205980 92150 206020 92350
rect 206090 92150 206410 92350
rect 206480 92150 206520 92350
rect 206590 92150 206910 92350
rect 206980 92150 207020 92350
rect 207090 92150 207410 92350
rect 207480 92150 207520 92350
rect 207590 92150 207910 92350
rect 207980 92150 208000 92350
rect 196000 92140 208000 92150
rect 196140 92090 196360 92140
rect 196140 92020 196150 92090
rect 196350 92020 196360 92090
rect 196140 91980 196360 92020
rect 196140 91910 196150 91980
rect 196350 91910 196360 91980
rect 196140 91860 196360 91910
rect 196640 92090 196860 92140
rect 196640 92020 196650 92090
rect 196850 92020 196860 92090
rect 196640 91980 196860 92020
rect 196640 91910 196650 91980
rect 196850 91910 196860 91980
rect 196640 91860 196860 91910
rect 197140 92090 197360 92140
rect 197140 92020 197150 92090
rect 197350 92020 197360 92090
rect 197140 91980 197360 92020
rect 197140 91910 197150 91980
rect 197350 91910 197360 91980
rect 197140 91860 197360 91910
rect 197640 92090 197860 92140
rect 197640 92020 197650 92090
rect 197850 92020 197860 92090
rect 197640 91980 197860 92020
rect 197640 91910 197650 91980
rect 197850 91910 197860 91980
rect 197640 91860 197860 91910
rect 198140 92090 198360 92140
rect 198140 92020 198150 92090
rect 198350 92020 198360 92090
rect 198140 91980 198360 92020
rect 198140 91910 198150 91980
rect 198350 91910 198360 91980
rect 198140 91860 198360 91910
rect 198640 92090 198860 92140
rect 198640 92020 198650 92090
rect 198850 92020 198860 92090
rect 198640 91980 198860 92020
rect 198640 91910 198650 91980
rect 198850 91910 198860 91980
rect 198640 91860 198860 91910
rect 199140 92090 199360 92140
rect 199140 92020 199150 92090
rect 199350 92020 199360 92090
rect 199140 91980 199360 92020
rect 199140 91910 199150 91980
rect 199350 91910 199360 91980
rect 199140 91860 199360 91910
rect 199640 92090 199860 92140
rect 199640 92020 199650 92090
rect 199850 92020 199860 92090
rect 199640 91980 199860 92020
rect 199640 91910 199650 91980
rect 199850 91910 199860 91980
rect 199640 91860 199860 91910
rect 200140 92090 200360 92140
rect 200140 92020 200150 92090
rect 200350 92020 200360 92090
rect 200140 91980 200360 92020
rect 200140 91910 200150 91980
rect 200350 91910 200360 91980
rect 200140 91860 200360 91910
rect 200640 92090 200860 92140
rect 200640 92020 200650 92090
rect 200850 92020 200860 92090
rect 200640 91980 200860 92020
rect 200640 91910 200650 91980
rect 200850 91910 200860 91980
rect 200640 91860 200860 91910
rect 201140 92090 201360 92140
rect 201140 92020 201150 92090
rect 201350 92020 201360 92090
rect 201140 91980 201360 92020
rect 201140 91910 201150 91980
rect 201350 91910 201360 91980
rect 201140 91860 201360 91910
rect 201640 92090 201860 92140
rect 201640 92020 201650 92090
rect 201850 92020 201860 92090
rect 201640 91980 201860 92020
rect 201640 91910 201650 91980
rect 201850 91910 201860 91980
rect 201640 91860 201860 91910
rect 202140 92090 202360 92140
rect 202140 92020 202150 92090
rect 202350 92020 202360 92090
rect 202140 91980 202360 92020
rect 202140 91910 202150 91980
rect 202350 91910 202360 91980
rect 202140 91860 202360 91910
rect 202640 92090 202860 92140
rect 202640 92020 202650 92090
rect 202850 92020 202860 92090
rect 202640 91980 202860 92020
rect 202640 91910 202650 91980
rect 202850 91910 202860 91980
rect 202640 91860 202860 91910
rect 203140 92090 203360 92140
rect 203140 92020 203150 92090
rect 203350 92020 203360 92090
rect 203140 91980 203360 92020
rect 203140 91910 203150 91980
rect 203350 91910 203360 91980
rect 203140 91860 203360 91910
rect 203640 92090 203860 92140
rect 203640 92020 203650 92090
rect 203850 92020 203860 92090
rect 203640 91980 203860 92020
rect 203640 91910 203650 91980
rect 203850 91910 203860 91980
rect 203640 91860 203860 91910
rect 204140 92090 204360 92140
rect 204140 92020 204150 92090
rect 204350 92020 204360 92090
rect 204140 91980 204360 92020
rect 204140 91910 204150 91980
rect 204350 91910 204360 91980
rect 204140 91860 204360 91910
rect 204640 92090 204860 92140
rect 204640 92020 204650 92090
rect 204850 92020 204860 92090
rect 204640 91980 204860 92020
rect 204640 91910 204650 91980
rect 204850 91910 204860 91980
rect 204640 91860 204860 91910
rect 205140 92090 205360 92140
rect 205140 92020 205150 92090
rect 205350 92020 205360 92090
rect 205140 91980 205360 92020
rect 205140 91910 205150 91980
rect 205350 91910 205360 91980
rect 205140 91860 205360 91910
rect 205640 92090 205860 92140
rect 205640 92020 205650 92090
rect 205850 92020 205860 92090
rect 205640 91980 205860 92020
rect 205640 91910 205650 91980
rect 205850 91910 205860 91980
rect 205640 91860 205860 91910
rect 206140 92090 206360 92140
rect 206140 92020 206150 92090
rect 206350 92020 206360 92090
rect 206140 91980 206360 92020
rect 206140 91910 206150 91980
rect 206350 91910 206360 91980
rect 206140 91860 206360 91910
rect 206640 92090 206860 92140
rect 206640 92020 206650 92090
rect 206850 92020 206860 92090
rect 206640 91980 206860 92020
rect 206640 91910 206650 91980
rect 206850 91910 206860 91980
rect 206640 91860 206860 91910
rect 207140 92090 207360 92140
rect 207140 92020 207150 92090
rect 207350 92020 207360 92090
rect 207140 91980 207360 92020
rect 207140 91910 207150 91980
rect 207350 91910 207360 91980
rect 207140 91860 207360 91910
rect 207640 92090 207860 92140
rect 207640 92020 207650 92090
rect 207850 92020 207860 92090
rect 207640 91980 207860 92020
rect 207640 91910 207650 91980
rect 207850 91910 207860 91980
rect 207640 91860 207860 91910
rect 196000 91850 208000 91860
rect 196000 91650 196020 91850
rect 196090 91650 196410 91850
rect 196480 91650 196520 91850
rect 196590 91650 196910 91850
rect 196980 91650 197020 91850
rect 197090 91650 197410 91850
rect 197480 91650 197520 91850
rect 197590 91650 197910 91850
rect 197980 91650 198020 91850
rect 198090 91650 198410 91850
rect 198480 91650 198520 91850
rect 198590 91650 198910 91850
rect 198980 91650 199020 91850
rect 199090 91650 199410 91850
rect 199480 91650 199520 91850
rect 199590 91650 199910 91850
rect 199980 91650 200020 91850
rect 200090 91650 200410 91850
rect 200480 91650 200520 91850
rect 200590 91650 200910 91850
rect 200980 91650 201020 91850
rect 201090 91650 201410 91850
rect 201480 91650 201520 91850
rect 201590 91650 201910 91850
rect 201980 91650 202020 91850
rect 202090 91650 202410 91850
rect 202480 91650 202520 91850
rect 202590 91650 202910 91850
rect 202980 91650 203020 91850
rect 203090 91650 203410 91850
rect 203480 91650 203520 91850
rect 203590 91650 203910 91850
rect 203980 91650 204020 91850
rect 204090 91650 204410 91850
rect 204480 91650 204520 91850
rect 204590 91650 204910 91850
rect 204980 91650 205020 91850
rect 205090 91650 205410 91850
rect 205480 91650 205520 91850
rect 205590 91650 205910 91850
rect 205980 91650 206020 91850
rect 206090 91650 206410 91850
rect 206480 91650 206520 91850
rect 206590 91650 206910 91850
rect 206980 91650 207020 91850
rect 207090 91650 207410 91850
rect 207480 91650 207520 91850
rect 207590 91650 207910 91850
rect 207980 91650 208000 91850
rect 196000 91640 208000 91650
rect 196140 91590 196360 91640
rect 196140 91520 196150 91590
rect 196350 91520 196360 91590
rect 196140 91480 196360 91520
rect 196140 91410 196150 91480
rect 196350 91410 196360 91480
rect 196140 91360 196360 91410
rect 196640 91590 196860 91640
rect 196640 91520 196650 91590
rect 196850 91520 196860 91590
rect 196640 91480 196860 91520
rect 196640 91410 196650 91480
rect 196850 91410 196860 91480
rect 196640 91360 196860 91410
rect 197140 91590 197360 91640
rect 197140 91520 197150 91590
rect 197350 91520 197360 91590
rect 197140 91480 197360 91520
rect 197140 91410 197150 91480
rect 197350 91410 197360 91480
rect 197140 91360 197360 91410
rect 197640 91590 197860 91640
rect 197640 91520 197650 91590
rect 197850 91520 197860 91590
rect 197640 91480 197860 91520
rect 197640 91410 197650 91480
rect 197850 91410 197860 91480
rect 197640 91360 197860 91410
rect 198140 91590 198360 91640
rect 198140 91520 198150 91590
rect 198350 91520 198360 91590
rect 198140 91480 198360 91520
rect 198140 91410 198150 91480
rect 198350 91410 198360 91480
rect 198140 91360 198360 91410
rect 198640 91590 198860 91640
rect 198640 91520 198650 91590
rect 198850 91520 198860 91590
rect 198640 91480 198860 91520
rect 198640 91410 198650 91480
rect 198850 91410 198860 91480
rect 198640 91360 198860 91410
rect 199140 91590 199360 91640
rect 199140 91520 199150 91590
rect 199350 91520 199360 91590
rect 199140 91480 199360 91520
rect 199140 91410 199150 91480
rect 199350 91410 199360 91480
rect 199140 91360 199360 91410
rect 199640 91590 199860 91640
rect 199640 91520 199650 91590
rect 199850 91520 199860 91590
rect 199640 91480 199860 91520
rect 199640 91410 199650 91480
rect 199850 91410 199860 91480
rect 199640 91360 199860 91410
rect 200140 91590 200360 91640
rect 200140 91520 200150 91590
rect 200350 91520 200360 91590
rect 200140 91480 200360 91520
rect 200140 91410 200150 91480
rect 200350 91410 200360 91480
rect 200140 91360 200360 91410
rect 200640 91590 200860 91640
rect 200640 91520 200650 91590
rect 200850 91520 200860 91590
rect 200640 91480 200860 91520
rect 200640 91410 200650 91480
rect 200850 91410 200860 91480
rect 200640 91360 200860 91410
rect 201140 91590 201360 91640
rect 201140 91520 201150 91590
rect 201350 91520 201360 91590
rect 201140 91480 201360 91520
rect 201140 91410 201150 91480
rect 201350 91410 201360 91480
rect 201140 91360 201360 91410
rect 201640 91590 201860 91640
rect 201640 91520 201650 91590
rect 201850 91520 201860 91590
rect 201640 91480 201860 91520
rect 201640 91410 201650 91480
rect 201850 91410 201860 91480
rect 201640 91360 201860 91410
rect 202140 91590 202360 91640
rect 202140 91520 202150 91590
rect 202350 91520 202360 91590
rect 202140 91480 202360 91520
rect 202140 91410 202150 91480
rect 202350 91410 202360 91480
rect 202140 91360 202360 91410
rect 202640 91590 202860 91640
rect 202640 91520 202650 91590
rect 202850 91520 202860 91590
rect 202640 91480 202860 91520
rect 202640 91410 202650 91480
rect 202850 91410 202860 91480
rect 202640 91360 202860 91410
rect 203140 91590 203360 91640
rect 203140 91520 203150 91590
rect 203350 91520 203360 91590
rect 203140 91480 203360 91520
rect 203140 91410 203150 91480
rect 203350 91410 203360 91480
rect 203140 91360 203360 91410
rect 203640 91590 203860 91640
rect 203640 91520 203650 91590
rect 203850 91520 203860 91590
rect 203640 91480 203860 91520
rect 203640 91410 203650 91480
rect 203850 91410 203860 91480
rect 203640 91360 203860 91410
rect 204140 91590 204360 91640
rect 204140 91520 204150 91590
rect 204350 91520 204360 91590
rect 204140 91480 204360 91520
rect 204140 91410 204150 91480
rect 204350 91410 204360 91480
rect 204140 91360 204360 91410
rect 204640 91590 204860 91640
rect 204640 91520 204650 91590
rect 204850 91520 204860 91590
rect 204640 91480 204860 91520
rect 204640 91410 204650 91480
rect 204850 91410 204860 91480
rect 204640 91360 204860 91410
rect 205140 91590 205360 91640
rect 205140 91520 205150 91590
rect 205350 91520 205360 91590
rect 205140 91480 205360 91520
rect 205140 91410 205150 91480
rect 205350 91410 205360 91480
rect 205140 91360 205360 91410
rect 205640 91590 205860 91640
rect 205640 91520 205650 91590
rect 205850 91520 205860 91590
rect 205640 91480 205860 91520
rect 205640 91410 205650 91480
rect 205850 91410 205860 91480
rect 205640 91360 205860 91410
rect 206140 91590 206360 91640
rect 206140 91520 206150 91590
rect 206350 91520 206360 91590
rect 206140 91480 206360 91520
rect 206140 91410 206150 91480
rect 206350 91410 206360 91480
rect 206140 91360 206360 91410
rect 206640 91590 206860 91640
rect 206640 91520 206650 91590
rect 206850 91520 206860 91590
rect 206640 91480 206860 91520
rect 206640 91410 206650 91480
rect 206850 91410 206860 91480
rect 206640 91360 206860 91410
rect 207140 91590 207360 91640
rect 207140 91520 207150 91590
rect 207350 91520 207360 91590
rect 207140 91480 207360 91520
rect 207140 91410 207150 91480
rect 207350 91410 207360 91480
rect 207140 91360 207360 91410
rect 207640 91590 207860 91640
rect 207640 91520 207650 91590
rect 207850 91520 207860 91590
rect 207640 91480 207860 91520
rect 207640 91410 207650 91480
rect 207850 91410 207860 91480
rect 207640 91360 207860 91410
rect 196000 91350 208000 91360
rect 196000 91150 196020 91350
rect 196090 91150 196410 91350
rect 196480 91150 196520 91350
rect 196590 91150 196910 91350
rect 196980 91150 197020 91350
rect 197090 91150 197410 91350
rect 197480 91150 197520 91350
rect 197590 91150 197910 91350
rect 197980 91150 198020 91350
rect 198090 91150 198410 91350
rect 198480 91150 198520 91350
rect 198590 91150 198910 91350
rect 198980 91150 199020 91350
rect 199090 91150 199410 91350
rect 199480 91150 199520 91350
rect 199590 91150 199910 91350
rect 199980 91150 200020 91350
rect 200090 91150 200410 91350
rect 200480 91150 200520 91350
rect 200590 91150 200910 91350
rect 200980 91150 201020 91350
rect 201090 91150 201410 91350
rect 201480 91150 201520 91350
rect 201590 91150 201910 91350
rect 201980 91150 202020 91350
rect 202090 91150 202410 91350
rect 202480 91150 202520 91350
rect 202590 91150 202910 91350
rect 202980 91150 203020 91350
rect 203090 91150 203410 91350
rect 203480 91150 203520 91350
rect 203590 91150 203910 91350
rect 203980 91150 204020 91350
rect 204090 91150 204410 91350
rect 204480 91150 204520 91350
rect 204590 91150 204910 91350
rect 204980 91150 205020 91350
rect 205090 91150 205410 91350
rect 205480 91150 205520 91350
rect 205590 91150 205910 91350
rect 205980 91150 206020 91350
rect 206090 91150 206410 91350
rect 206480 91150 206520 91350
rect 206590 91150 206910 91350
rect 206980 91150 207020 91350
rect 207090 91150 207410 91350
rect 207480 91150 207520 91350
rect 207590 91150 207910 91350
rect 207980 91150 208000 91350
rect 196000 91140 208000 91150
rect 196140 91090 196360 91140
rect 196140 91020 196150 91090
rect 196350 91020 196360 91090
rect 196140 90980 196360 91020
rect 196140 90910 196150 90980
rect 196350 90910 196360 90980
rect 196140 90860 196360 90910
rect 196640 91090 196860 91140
rect 196640 91020 196650 91090
rect 196850 91020 196860 91090
rect 196640 90980 196860 91020
rect 196640 90910 196650 90980
rect 196850 90910 196860 90980
rect 196640 90860 196860 90910
rect 197140 91090 197360 91140
rect 197140 91020 197150 91090
rect 197350 91020 197360 91090
rect 197140 90980 197360 91020
rect 197140 90910 197150 90980
rect 197350 90910 197360 90980
rect 197140 90860 197360 90910
rect 197640 91090 197860 91140
rect 197640 91020 197650 91090
rect 197850 91020 197860 91090
rect 197640 90980 197860 91020
rect 197640 90910 197650 90980
rect 197850 90910 197860 90980
rect 197640 90860 197860 90910
rect 198140 91090 198360 91140
rect 198140 91020 198150 91090
rect 198350 91020 198360 91090
rect 198140 90980 198360 91020
rect 198140 90910 198150 90980
rect 198350 90910 198360 90980
rect 198140 90860 198360 90910
rect 198640 91090 198860 91140
rect 198640 91020 198650 91090
rect 198850 91020 198860 91090
rect 198640 90980 198860 91020
rect 198640 90910 198650 90980
rect 198850 90910 198860 90980
rect 198640 90860 198860 90910
rect 199140 91090 199360 91140
rect 199140 91020 199150 91090
rect 199350 91020 199360 91090
rect 199140 90980 199360 91020
rect 199140 90910 199150 90980
rect 199350 90910 199360 90980
rect 199140 90860 199360 90910
rect 199640 91090 199860 91140
rect 199640 91020 199650 91090
rect 199850 91020 199860 91090
rect 199640 90980 199860 91020
rect 199640 90910 199650 90980
rect 199850 90910 199860 90980
rect 199640 90860 199860 90910
rect 200140 91090 200360 91140
rect 200140 91020 200150 91090
rect 200350 91020 200360 91090
rect 200140 90980 200360 91020
rect 200140 90910 200150 90980
rect 200350 90910 200360 90980
rect 200140 90860 200360 90910
rect 200640 91090 200860 91140
rect 200640 91020 200650 91090
rect 200850 91020 200860 91090
rect 200640 90980 200860 91020
rect 200640 90910 200650 90980
rect 200850 90910 200860 90980
rect 200640 90860 200860 90910
rect 201140 91090 201360 91140
rect 201140 91020 201150 91090
rect 201350 91020 201360 91090
rect 201140 90980 201360 91020
rect 201140 90910 201150 90980
rect 201350 90910 201360 90980
rect 201140 90860 201360 90910
rect 201640 91090 201860 91140
rect 201640 91020 201650 91090
rect 201850 91020 201860 91090
rect 201640 90980 201860 91020
rect 201640 90910 201650 90980
rect 201850 90910 201860 90980
rect 201640 90860 201860 90910
rect 202140 91090 202360 91140
rect 202140 91020 202150 91090
rect 202350 91020 202360 91090
rect 202140 90980 202360 91020
rect 202140 90910 202150 90980
rect 202350 90910 202360 90980
rect 202140 90860 202360 90910
rect 202640 91090 202860 91140
rect 202640 91020 202650 91090
rect 202850 91020 202860 91090
rect 202640 90980 202860 91020
rect 202640 90910 202650 90980
rect 202850 90910 202860 90980
rect 202640 90860 202860 90910
rect 203140 91090 203360 91140
rect 203140 91020 203150 91090
rect 203350 91020 203360 91090
rect 203140 90980 203360 91020
rect 203140 90910 203150 90980
rect 203350 90910 203360 90980
rect 203140 90860 203360 90910
rect 203640 91090 203860 91140
rect 203640 91020 203650 91090
rect 203850 91020 203860 91090
rect 203640 90980 203860 91020
rect 203640 90910 203650 90980
rect 203850 90910 203860 90980
rect 203640 90860 203860 90910
rect 204140 91090 204360 91140
rect 204140 91020 204150 91090
rect 204350 91020 204360 91090
rect 204140 90980 204360 91020
rect 204140 90910 204150 90980
rect 204350 90910 204360 90980
rect 204140 90860 204360 90910
rect 204640 91090 204860 91140
rect 204640 91020 204650 91090
rect 204850 91020 204860 91090
rect 204640 90980 204860 91020
rect 204640 90910 204650 90980
rect 204850 90910 204860 90980
rect 204640 90860 204860 90910
rect 205140 91090 205360 91140
rect 205140 91020 205150 91090
rect 205350 91020 205360 91090
rect 205140 90980 205360 91020
rect 205140 90910 205150 90980
rect 205350 90910 205360 90980
rect 205140 90860 205360 90910
rect 205640 91090 205860 91140
rect 205640 91020 205650 91090
rect 205850 91020 205860 91090
rect 205640 90980 205860 91020
rect 205640 90910 205650 90980
rect 205850 90910 205860 90980
rect 205640 90860 205860 90910
rect 206140 91090 206360 91140
rect 206140 91020 206150 91090
rect 206350 91020 206360 91090
rect 206140 90980 206360 91020
rect 206140 90910 206150 90980
rect 206350 90910 206360 90980
rect 206140 90860 206360 90910
rect 206640 91090 206860 91140
rect 206640 91020 206650 91090
rect 206850 91020 206860 91090
rect 206640 90980 206860 91020
rect 206640 90910 206650 90980
rect 206850 90910 206860 90980
rect 206640 90860 206860 90910
rect 207140 91090 207360 91140
rect 207140 91020 207150 91090
rect 207350 91020 207360 91090
rect 207140 90980 207360 91020
rect 207140 90910 207150 90980
rect 207350 90910 207360 90980
rect 207140 90860 207360 90910
rect 207640 91090 207860 91140
rect 207640 91020 207650 91090
rect 207850 91020 207860 91090
rect 207640 90980 207860 91020
rect 207640 90910 207650 90980
rect 207850 90910 207860 90980
rect 207640 90860 207860 90910
rect 196000 90850 208000 90860
rect 196000 90650 196020 90850
rect 196090 90650 196410 90850
rect 196480 90650 196520 90850
rect 196590 90650 196910 90850
rect 196980 90650 197020 90850
rect 197090 90650 197410 90850
rect 197480 90650 197520 90850
rect 197590 90650 197910 90850
rect 197980 90650 198020 90850
rect 198090 90650 198410 90850
rect 198480 90650 198520 90850
rect 198590 90650 198910 90850
rect 198980 90650 199020 90850
rect 199090 90650 199410 90850
rect 199480 90650 199520 90850
rect 199590 90650 199910 90850
rect 199980 90650 200020 90850
rect 200090 90650 200410 90850
rect 200480 90650 200520 90850
rect 200590 90650 200910 90850
rect 200980 90650 201020 90850
rect 201090 90650 201410 90850
rect 201480 90650 201520 90850
rect 201590 90650 201910 90850
rect 201980 90650 202020 90850
rect 202090 90650 202410 90850
rect 202480 90650 202520 90850
rect 202590 90650 202910 90850
rect 202980 90650 203020 90850
rect 203090 90650 203410 90850
rect 203480 90650 203520 90850
rect 203590 90650 203910 90850
rect 203980 90650 204020 90850
rect 204090 90650 204410 90850
rect 204480 90650 204520 90850
rect 204590 90650 204910 90850
rect 204980 90650 205020 90850
rect 205090 90650 205410 90850
rect 205480 90650 205520 90850
rect 205590 90650 205910 90850
rect 205980 90650 206020 90850
rect 206090 90650 206410 90850
rect 206480 90650 206520 90850
rect 206590 90650 206910 90850
rect 206980 90650 207020 90850
rect 207090 90650 207410 90850
rect 207480 90650 207520 90850
rect 207590 90650 207910 90850
rect 207980 90650 208000 90850
rect 196000 90640 208000 90650
rect 196140 90590 196360 90640
rect 196140 90520 196150 90590
rect 196350 90520 196360 90590
rect 196140 90480 196360 90520
rect 196140 90410 196150 90480
rect 196350 90410 196360 90480
rect 196140 90360 196360 90410
rect 196640 90590 196860 90640
rect 196640 90520 196650 90590
rect 196850 90520 196860 90590
rect 196640 90480 196860 90520
rect 196640 90410 196650 90480
rect 196850 90410 196860 90480
rect 196640 90360 196860 90410
rect 197140 90590 197360 90640
rect 197140 90520 197150 90590
rect 197350 90520 197360 90590
rect 197140 90480 197360 90520
rect 197140 90410 197150 90480
rect 197350 90410 197360 90480
rect 197140 90360 197360 90410
rect 197640 90590 197860 90640
rect 197640 90520 197650 90590
rect 197850 90520 197860 90590
rect 197640 90480 197860 90520
rect 197640 90410 197650 90480
rect 197850 90410 197860 90480
rect 197640 90360 197860 90410
rect 198140 90590 198360 90640
rect 198140 90520 198150 90590
rect 198350 90520 198360 90590
rect 198140 90480 198360 90520
rect 198140 90410 198150 90480
rect 198350 90410 198360 90480
rect 198140 90360 198360 90410
rect 198640 90590 198860 90640
rect 198640 90520 198650 90590
rect 198850 90520 198860 90590
rect 198640 90480 198860 90520
rect 198640 90410 198650 90480
rect 198850 90410 198860 90480
rect 198640 90360 198860 90410
rect 199140 90590 199360 90640
rect 199140 90520 199150 90590
rect 199350 90520 199360 90590
rect 199140 90480 199360 90520
rect 199140 90410 199150 90480
rect 199350 90410 199360 90480
rect 199140 90360 199360 90410
rect 199640 90590 199860 90640
rect 199640 90520 199650 90590
rect 199850 90520 199860 90590
rect 199640 90480 199860 90520
rect 199640 90410 199650 90480
rect 199850 90410 199860 90480
rect 199640 90360 199860 90410
rect 200140 90590 200360 90640
rect 200140 90520 200150 90590
rect 200350 90520 200360 90590
rect 200140 90480 200360 90520
rect 200140 90410 200150 90480
rect 200350 90410 200360 90480
rect 200140 90360 200360 90410
rect 200640 90590 200860 90640
rect 200640 90520 200650 90590
rect 200850 90520 200860 90590
rect 200640 90480 200860 90520
rect 200640 90410 200650 90480
rect 200850 90410 200860 90480
rect 200640 90360 200860 90410
rect 201140 90590 201360 90640
rect 201140 90520 201150 90590
rect 201350 90520 201360 90590
rect 201140 90480 201360 90520
rect 201140 90410 201150 90480
rect 201350 90410 201360 90480
rect 201140 90360 201360 90410
rect 201640 90590 201860 90640
rect 201640 90520 201650 90590
rect 201850 90520 201860 90590
rect 201640 90480 201860 90520
rect 201640 90410 201650 90480
rect 201850 90410 201860 90480
rect 201640 90360 201860 90410
rect 202140 90590 202360 90640
rect 202140 90520 202150 90590
rect 202350 90520 202360 90590
rect 202140 90480 202360 90520
rect 202140 90410 202150 90480
rect 202350 90410 202360 90480
rect 202140 90360 202360 90410
rect 202640 90590 202860 90640
rect 202640 90520 202650 90590
rect 202850 90520 202860 90590
rect 202640 90480 202860 90520
rect 202640 90410 202650 90480
rect 202850 90410 202860 90480
rect 202640 90360 202860 90410
rect 203140 90590 203360 90640
rect 203140 90520 203150 90590
rect 203350 90520 203360 90590
rect 203140 90480 203360 90520
rect 203140 90410 203150 90480
rect 203350 90410 203360 90480
rect 203140 90360 203360 90410
rect 203640 90590 203860 90640
rect 203640 90520 203650 90590
rect 203850 90520 203860 90590
rect 203640 90480 203860 90520
rect 203640 90410 203650 90480
rect 203850 90410 203860 90480
rect 203640 90360 203860 90410
rect 204140 90590 204360 90640
rect 204140 90520 204150 90590
rect 204350 90520 204360 90590
rect 204140 90480 204360 90520
rect 204140 90410 204150 90480
rect 204350 90410 204360 90480
rect 204140 90360 204360 90410
rect 204640 90590 204860 90640
rect 204640 90520 204650 90590
rect 204850 90520 204860 90590
rect 204640 90480 204860 90520
rect 204640 90410 204650 90480
rect 204850 90410 204860 90480
rect 204640 90360 204860 90410
rect 205140 90590 205360 90640
rect 205140 90520 205150 90590
rect 205350 90520 205360 90590
rect 205140 90480 205360 90520
rect 205140 90410 205150 90480
rect 205350 90410 205360 90480
rect 205140 90360 205360 90410
rect 205640 90590 205860 90640
rect 205640 90520 205650 90590
rect 205850 90520 205860 90590
rect 205640 90480 205860 90520
rect 205640 90410 205650 90480
rect 205850 90410 205860 90480
rect 205640 90360 205860 90410
rect 206140 90590 206360 90640
rect 206140 90520 206150 90590
rect 206350 90520 206360 90590
rect 206140 90480 206360 90520
rect 206140 90410 206150 90480
rect 206350 90410 206360 90480
rect 206140 90360 206360 90410
rect 206640 90590 206860 90640
rect 206640 90520 206650 90590
rect 206850 90520 206860 90590
rect 206640 90480 206860 90520
rect 206640 90410 206650 90480
rect 206850 90410 206860 90480
rect 206640 90360 206860 90410
rect 207140 90590 207360 90640
rect 207140 90520 207150 90590
rect 207350 90520 207360 90590
rect 207140 90480 207360 90520
rect 207140 90410 207150 90480
rect 207350 90410 207360 90480
rect 207140 90360 207360 90410
rect 207640 90590 207860 90640
rect 207640 90520 207650 90590
rect 207850 90520 207860 90590
rect 207640 90480 207860 90520
rect 207640 90410 207650 90480
rect 207850 90410 207860 90480
rect 207640 90360 207860 90410
rect 196000 90350 208000 90360
rect 196000 90150 196020 90350
rect 196090 90150 196410 90350
rect 196480 90150 196520 90350
rect 196590 90150 196910 90350
rect 196980 90150 197020 90350
rect 197090 90150 197410 90350
rect 197480 90150 197520 90350
rect 197590 90150 197910 90350
rect 197980 90150 198020 90350
rect 198090 90150 198410 90350
rect 198480 90150 198520 90350
rect 198590 90150 198910 90350
rect 198980 90150 199020 90350
rect 199090 90150 199410 90350
rect 199480 90150 199520 90350
rect 199590 90150 199910 90350
rect 199980 90150 200020 90350
rect 200090 90150 200410 90350
rect 200480 90150 200520 90350
rect 200590 90150 200910 90350
rect 200980 90150 201020 90350
rect 201090 90150 201410 90350
rect 201480 90150 201520 90350
rect 201590 90150 201910 90350
rect 201980 90150 202020 90350
rect 202090 90150 202410 90350
rect 202480 90150 202520 90350
rect 202590 90150 202910 90350
rect 202980 90150 203020 90350
rect 203090 90150 203410 90350
rect 203480 90150 203520 90350
rect 203590 90150 203910 90350
rect 203980 90150 204020 90350
rect 204090 90150 204410 90350
rect 204480 90150 204520 90350
rect 204590 90150 204910 90350
rect 204980 90150 205020 90350
rect 205090 90150 205410 90350
rect 205480 90150 205520 90350
rect 205590 90150 205910 90350
rect 205980 90150 206020 90350
rect 206090 90150 206410 90350
rect 206480 90150 206520 90350
rect 206590 90150 206910 90350
rect 206980 90150 207020 90350
rect 207090 90150 207410 90350
rect 207480 90150 207520 90350
rect 207590 90150 207910 90350
rect 207980 90150 208000 90350
rect 196000 90140 208000 90150
rect 196140 90090 196360 90140
rect 196140 90020 196150 90090
rect 196350 90020 196360 90090
rect 196140 89980 196360 90020
rect 196140 89910 196150 89980
rect 196350 89910 196360 89980
rect 196140 89860 196360 89910
rect 196640 90090 196860 90140
rect 196640 90020 196650 90090
rect 196850 90020 196860 90090
rect 196640 89980 196860 90020
rect 196640 89910 196650 89980
rect 196850 89910 196860 89980
rect 196640 89860 196860 89910
rect 197140 90090 197360 90140
rect 197140 90020 197150 90090
rect 197350 90020 197360 90090
rect 197140 89980 197360 90020
rect 197140 89910 197150 89980
rect 197350 89910 197360 89980
rect 197140 89860 197360 89910
rect 197640 90090 197860 90140
rect 197640 90020 197650 90090
rect 197850 90020 197860 90090
rect 197640 89980 197860 90020
rect 197640 89910 197650 89980
rect 197850 89910 197860 89980
rect 197640 89860 197860 89910
rect 198140 90090 198360 90140
rect 198140 90020 198150 90090
rect 198350 90020 198360 90090
rect 198140 89980 198360 90020
rect 198140 89910 198150 89980
rect 198350 89910 198360 89980
rect 198140 89860 198360 89910
rect 198640 90090 198860 90140
rect 198640 90020 198650 90090
rect 198850 90020 198860 90090
rect 198640 89980 198860 90020
rect 198640 89910 198650 89980
rect 198850 89910 198860 89980
rect 198640 89860 198860 89910
rect 199140 90090 199360 90140
rect 199140 90020 199150 90090
rect 199350 90020 199360 90090
rect 199140 89980 199360 90020
rect 199140 89910 199150 89980
rect 199350 89910 199360 89980
rect 199140 89860 199360 89910
rect 199640 90090 199860 90140
rect 199640 90020 199650 90090
rect 199850 90020 199860 90090
rect 199640 89980 199860 90020
rect 199640 89910 199650 89980
rect 199850 89910 199860 89980
rect 199640 89860 199860 89910
rect 200140 90090 200360 90140
rect 200140 90020 200150 90090
rect 200350 90020 200360 90090
rect 200140 89980 200360 90020
rect 200140 89910 200150 89980
rect 200350 89910 200360 89980
rect 200140 89860 200360 89910
rect 200640 90090 200860 90140
rect 200640 90020 200650 90090
rect 200850 90020 200860 90090
rect 200640 89980 200860 90020
rect 200640 89910 200650 89980
rect 200850 89910 200860 89980
rect 200640 89860 200860 89910
rect 201140 90090 201360 90140
rect 201140 90020 201150 90090
rect 201350 90020 201360 90090
rect 201140 89980 201360 90020
rect 201140 89910 201150 89980
rect 201350 89910 201360 89980
rect 201140 89860 201360 89910
rect 201640 90090 201860 90140
rect 201640 90020 201650 90090
rect 201850 90020 201860 90090
rect 201640 89980 201860 90020
rect 201640 89910 201650 89980
rect 201850 89910 201860 89980
rect 201640 89860 201860 89910
rect 202140 90090 202360 90140
rect 202140 90020 202150 90090
rect 202350 90020 202360 90090
rect 202140 89980 202360 90020
rect 202140 89910 202150 89980
rect 202350 89910 202360 89980
rect 202140 89860 202360 89910
rect 202640 90090 202860 90140
rect 202640 90020 202650 90090
rect 202850 90020 202860 90090
rect 202640 89980 202860 90020
rect 202640 89910 202650 89980
rect 202850 89910 202860 89980
rect 202640 89860 202860 89910
rect 203140 90090 203360 90140
rect 203140 90020 203150 90090
rect 203350 90020 203360 90090
rect 203140 89980 203360 90020
rect 203140 89910 203150 89980
rect 203350 89910 203360 89980
rect 203140 89860 203360 89910
rect 203640 90090 203860 90140
rect 203640 90020 203650 90090
rect 203850 90020 203860 90090
rect 203640 89980 203860 90020
rect 203640 89910 203650 89980
rect 203850 89910 203860 89980
rect 203640 89860 203860 89910
rect 204140 90090 204360 90140
rect 204140 90020 204150 90090
rect 204350 90020 204360 90090
rect 204140 89980 204360 90020
rect 204140 89910 204150 89980
rect 204350 89910 204360 89980
rect 204140 89860 204360 89910
rect 204640 90090 204860 90140
rect 204640 90020 204650 90090
rect 204850 90020 204860 90090
rect 204640 89980 204860 90020
rect 204640 89910 204650 89980
rect 204850 89910 204860 89980
rect 204640 89860 204860 89910
rect 205140 90090 205360 90140
rect 205140 90020 205150 90090
rect 205350 90020 205360 90090
rect 205140 89980 205360 90020
rect 205140 89910 205150 89980
rect 205350 89910 205360 89980
rect 205140 89860 205360 89910
rect 205640 90090 205860 90140
rect 205640 90020 205650 90090
rect 205850 90020 205860 90090
rect 205640 89980 205860 90020
rect 205640 89910 205650 89980
rect 205850 89910 205860 89980
rect 205640 89860 205860 89910
rect 206140 90090 206360 90140
rect 206140 90020 206150 90090
rect 206350 90020 206360 90090
rect 206140 89980 206360 90020
rect 206140 89910 206150 89980
rect 206350 89910 206360 89980
rect 206140 89860 206360 89910
rect 206640 90090 206860 90140
rect 206640 90020 206650 90090
rect 206850 90020 206860 90090
rect 206640 89980 206860 90020
rect 206640 89910 206650 89980
rect 206850 89910 206860 89980
rect 206640 89860 206860 89910
rect 207140 90090 207360 90140
rect 207140 90020 207150 90090
rect 207350 90020 207360 90090
rect 207140 89980 207360 90020
rect 207140 89910 207150 89980
rect 207350 89910 207360 89980
rect 207140 89860 207360 89910
rect 207640 90090 207860 90140
rect 207640 90020 207650 90090
rect 207850 90020 207860 90090
rect 207640 89980 207860 90020
rect 207640 89910 207650 89980
rect 207850 89910 207860 89980
rect 207640 89860 207860 89910
rect 196000 89850 208000 89860
rect 196000 89650 196020 89850
rect 196090 89650 196410 89850
rect 196480 89650 196520 89850
rect 196590 89650 196910 89850
rect 196980 89650 197020 89850
rect 197090 89650 197410 89850
rect 197480 89650 197520 89850
rect 197590 89650 197910 89850
rect 197980 89650 198020 89850
rect 198090 89650 198410 89850
rect 198480 89650 198520 89850
rect 198590 89650 198910 89850
rect 198980 89650 199020 89850
rect 199090 89650 199410 89850
rect 199480 89650 199520 89850
rect 199590 89650 199910 89850
rect 199980 89650 200020 89850
rect 200090 89650 200410 89850
rect 200480 89650 200520 89850
rect 200590 89650 200910 89850
rect 200980 89650 201020 89850
rect 201090 89650 201410 89850
rect 201480 89650 201520 89850
rect 201590 89650 201910 89850
rect 201980 89650 202020 89850
rect 202090 89650 202410 89850
rect 202480 89650 202520 89850
rect 202590 89650 202910 89850
rect 202980 89650 203020 89850
rect 203090 89650 203410 89850
rect 203480 89650 203520 89850
rect 203590 89650 203910 89850
rect 203980 89650 204020 89850
rect 204090 89650 204410 89850
rect 204480 89650 204520 89850
rect 204590 89650 204910 89850
rect 204980 89650 205020 89850
rect 205090 89650 205410 89850
rect 205480 89650 205520 89850
rect 205590 89650 205910 89850
rect 205980 89650 206020 89850
rect 206090 89650 206410 89850
rect 206480 89650 206520 89850
rect 206590 89650 206910 89850
rect 206980 89650 207020 89850
rect 207090 89650 207410 89850
rect 207480 89650 207520 89850
rect 207590 89650 207910 89850
rect 207980 89650 208000 89850
rect 196000 89640 208000 89650
rect 196140 89590 196360 89640
rect 196140 89520 196150 89590
rect 196350 89520 196360 89590
rect 196140 89480 196360 89520
rect 196140 89410 196150 89480
rect 196350 89410 196360 89480
rect 196140 89360 196360 89410
rect 196640 89590 196860 89640
rect 196640 89520 196650 89590
rect 196850 89520 196860 89590
rect 196640 89480 196860 89520
rect 196640 89410 196650 89480
rect 196850 89410 196860 89480
rect 196640 89360 196860 89410
rect 197140 89590 197360 89640
rect 197140 89520 197150 89590
rect 197350 89520 197360 89590
rect 197140 89480 197360 89520
rect 197140 89410 197150 89480
rect 197350 89410 197360 89480
rect 197140 89360 197360 89410
rect 197640 89590 197860 89640
rect 197640 89520 197650 89590
rect 197850 89520 197860 89590
rect 197640 89480 197860 89520
rect 197640 89410 197650 89480
rect 197850 89410 197860 89480
rect 197640 89360 197860 89410
rect 198140 89590 198360 89640
rect 198140 89520 198150 89590
rect 198350 89520 198360 89590
rect 198140 89480 198360 89520
rect 198140 89410 198150 89480
rect 198350 89410 198360 89480
rect 198140 89360 198360 89410
rect 198640 89590 198860 89640
rect 198640 89520 198650 89590
rect 198850 89520 198860 89590
rect 198640 89480 198860 89520
rect 198640 89410 198650 89480
rect 198850 89410 198860 89480
rect 198640 89360 198860 89410
rect 199140 89590 199360 89640
rect 199140 89520 199150 89590
rect 199350 89520 199360 89590
rect 199140 89480 199360 89520
rect 199140 89410 199150 89480
rect 199350 89410 199360 89480
rect 199140 89360 199360 89410
rect 199640 89590 199860 89640
rect 199640 89520 199650 89590
rect 199850 89520 199860 89590
rect 199640 89480 199860 89520
rect 199640 89410 199650 89480
rect 199850 89410 199860 89480
rect 199640 89360 199860 89410
rect 200140 89590 200360 89640
rect 200140 89520 200150 89590
rect 200350 89520 200360 89590
rect 200140 89480 200360 89520
rect 200140 89410 200150 89480
rect 200350 89410 200360 89480
rect 200140 89360 200360 89410
rect 200640 89590 200860 89640
rect 200640 89520 200650 89590
rect 200850 89520 200860 89590
rect 200640 89480 200860 89520
rect 200640 89410 200650 89480
rect 200850 89410 200860 89480
rect 200640 89360 200860 89410
rect 201140 89590 201360 89640
rect 201140 89520 201150 89590
rect 201350 89520 201360 89590
rect 201140 89480 201360 89520
rect 201140 89410 201150 89480
rect 201350 89410 201360 89480
rect 201140 89360 201360 89410
rect 201640 89590 201860 89640
rect 201640 89520 201650 89590
rect 201850 89520 201860 89590
rect 201640 89480 201860 89520
rect 201640 89410 201650 89480
rect 201850 89410 201860 89480
rect 201640 89360 201860 89410
rect 202140 89590 202360 89640
rect 202140 89520 202150 89590
rect 202350 89520 202360 89590
rect 202140 89480 202360 89520
rect 202140 89410 202150 89480
rect 202350 89410 202360 89480
rect 202140 89360 202360 89410
rect 202640 89590 202860 89640
rect 202640 89520 202650 89590
rect 202850 89520 202860 89590
rect 202640 89480 202860 89520
rect 202640 89410 202650 89480
rect 202850 89410 202860 89480
rect 202640 89360 202860 89410
rect 203140 89590 203360 89640
rect 203140 89520 203150 89590
rect 203350 89520 203360 89590
rect 203140 89480 203360 89520
rect 203140 89410 203150 89480
rect 203350 89410 203360 89480
rect 203140 89360 203360 89410
rect 203640 89590 203860 89640
rect 203640 89520 203650 89590
rect 203850 89520 203860 89590
rect 203640 89480 203860 89520
rect 203640 89410 203650 89480
rect 203850 89410 203860 89480
rect 203640 89360 203860 89410
rect 204140 89590 204360 89640
rect 204140 89520 204150 89590
rect 204350 89520 204360 89590
rect 204140 89480 204360 89520
rect 204140 89410 204150 89480
rect 204350 89410 204360 89480
rect 204140 89360 204360 89410
rect 204640 89590 204860 89640
rect 204640 89520 204650 89590
rect 204850 89520 204860 89590
rect 204640 89480 204860 89520
rect 204640 89410 204650 89480
rect 204850 89410 204860 89480
rect 204640 89360 204860 89410
rect 205140 89590 205360 89640
rect 205140 89520 205150 89590
rect 205350 89520 205360 89590
rect 205140 89480 205360 89520
rect 205140 89410 205150 89480
rect 205350 89410 205360 89480
rect 205140 89360 205360 89410
rect 205640 89590 205860 89640
rect 205640 89520 205650 89590
rect 205850 89520 205860 89590
rect 205640 89480 205860 89520
rect 205640 89410 205650 89480
rect 205850 89410 205860 89480
rect 205640 89360 205860 89410
rect 206140 89590 206360 89640
rect 206140 89520 206150 89590
rect 206350 89520 206360 89590
rect 206140 89480 206360 89520
rect 206140 89410 206150 89480
rect 206350 89410 206360 89480
rect 206140 89360 206360 89410
rect 206640 89590 206860 89640
rect 206640 89520 206650 89590
rect 206850 89520 206860 89590
rect 206640 89480 206860 89520
rect 206640 89410 206650 89480
rect 206850 89410 206860 89480
rect 206640 89360 206860 89410
rect 207140 89590 207360 89640
rect 207140 89520 207150 89590
rect 207350 89520 207360 89590
rect 207140 89480 207360 89520
rect 207140 89410 207150 89480
rect 207350 89410 207360 89480
rect 207140 89360 207360 89410
rect 207640 89590 207860 89640
rect 207640 89520 207650 89590
rect 207850 89520 207860 89590
rect 207640 89480 207860 89520
rect 207640 89410 207650 89480
rect 207850 89410 207860 89480
rect 207640 89360 207860 89410
rect 196000 89350 208000 89360
rect 196000 89150 196020 89350
rect 196090 89150 196410 89350
rect 196480 89150 196520 89350
rect 196590 89150 196910 89350
rect 196980 89150 197020 89350
rect 197090 89150 197410 89350
rect 197480 89150 197520 89350
rect 197590 89150 197910 89350
rect 197980 89150 198020 89350
rect 198090 89150 198410 89350
rect 198480 89150 198520 89350
rect 198590 89150 198910 89350
rect 198980 89150 199020 89350
rect 199090 89150 199410 89350
rect 199480 89150 199520 89350
rect 199590 89150 199910 89350
rect 199980 89150 200020 89350
rect 200090 89150 200410 89350
rect 200480 89150 200520 89350
rect 200590 89150 200910 89350
rect 200980 89150 201020 89350
rect 201090 89150 201410 89350
rect 201480 89150 201520 89350
rect 201590 89150 201910 89350
rect 201980 89150 202020 89350
rect 202090 89150 202410 89350
rect 202480 89150 202520 89350
rect 202590 89150 202910 89350
rect 202980 89150 203020 89350
rect 203090 89150 203410 89350
rect 203480 89150 203520 89350
rect 203590 89150 203910 89350
rect 203980 89150 204020 89350
rect 204090 89150 204410 89350
rect 204480 89150 204520 89350
rect 204590 89150 204910 89350
rect 204980 89150 205020 89350
rect 205090 89150 205410 89350
rect 205480 89150 205520 89350
rect 205590 89150 205910 89350
rect 205980 89150 206020 89350
rect 206090 89150 206410 89350
rect 206480 89150 206520 89350
rect 206590 89150 206910 89350
rect 206980 89150 207020 89350
rect 207090 89150 207410 89350
rect 207480 89150 207520 89350
rect 207590 89150 207910 89350
rect 207980 89150 208000 89350
rect 196000 89140 208000 89150
rect 196140 89090 196360 89140
rect 196140 89020 196150 89090
rect 196350 89020 196360 89090
rect 196140 88980 196360 89020
rect 196140 88910 196150 88980
rect 196350 88910 196360 88980
rect 196140 88860 196360 88910
rect 196640 89090 196860 89140
rect 196640 89020 196650 89090
rect 196850 89020 196860 89090
rect 196640 88980 196860 89020
rect 196640 88910 196650 88980
rect 196850 88910 196860 88980
rect 196640 88860 196860 88910
rect 197140 89090 197360 89140
rect 197140 89020 197150 89090
rect 197350 89020 197360 89090
rect 197140 88980 197360 89020
rect 197140 88910 197150 88980
rect 197350 88910 197360 88980
rect 197140 88860 197360 88910
rect 197640 89090 197860 89140
rect 197640 89020 197650 89090
rect 197850 89020 197860 89090
rect 197640 88980 197860 89020
rect 197640 88910 197650 88980
rect 197850 88910 197860 88980
rect 197640 88860 197860 88910
rect 198140 89090 198360 89140
rect 198140 89020 198150 89090
rect 198350 89020 198360 89090
rect 198140 88980 198360 89020
rect 198140 88910 198150 88980
rect 198350 88910 198360 88980
rect 198140 88860 198360 88910
rect 198640 89090 198860 89140
rect 198640 89020 198650 89090
rect 198850 89020 198860 89090
rect 198640 88980 198860 89020
rect 198640 88910 198650 88980
rect 198850 88910 198860 88980
rect 198640 88860 198860 88910
rect 199140 89090 199360 89140
rect 199140 89020 199150 89090
rect 199350 89020 199360 89090
rect 199140 88980 199360 89020
rect 199140 88910 199150 88980
rect 199350 88910 199360 88980
rect 199140 88860 199360 88910
rect 199640 89090 199860 89140
rect 199640 89020 199650 89090
rect 199850 89020 199860 89090
rect 199640 88980 199860 89020
rect 199640 88910 199650 88980
rect 199850 88910 199860 88980
rect 199640 88860 199860 88910
rect 200140 89090 200360 89140
rect 200140 89020 200150 89090
rect 200350 89020 200360 89090
rect 200140 88980 200360 89020
rect 200140 88910 200150 88980
rect 200350 88910 200360 88980
rect 200140 88860 200360 88910
rect 200640 89090 200860 89140
rect 200640 89020 200650 89090
rect 200850 89020 200860 89090
rect 200640 88980 200860 89020
rect 200640 88910 200650 88980
rect 200850 88910 200860 88980
rect 200640 88860 200860 88910
rect 201140 89090 201360 89140
rect 201140 89020 201150 89090
rect 201350 89020 201360 89090
rect 201140 88980 201360 89020
rect 201140 88910 201150 88980
rect 201350 88910 201360 88980
rect 201140 88860 201360 88910
rect 201640 89090 201860 89140
rect 201640 89020 201650 89090
rect 201850 89020 201860 89090
rect 201640 88980 201860 89020
rect 201640 88910 201650 88980
rect 201850 88910 201860 88980
rect 201640 88860 201860 88910
rect 202140 89090 202360 89140
rect 202140 89020 202150 89090
rect 202350 89020 202360 89090
rect 202140 88980 202360 89020
rect 202140 88910 202150 88980
rect 202350 88910 202360 88980
rect 202140 88860 202360 88910
rect 202640 89090 202860 89140
rect 202640 89020 202650 89090
rect 202850 89020 202860 89090
rect 202640 88980 202860 89020
rect 202640 88910 202650 88980
rect 202850 88910 202860 88980
rect 202640 88860 202860 88910
rect 203140 89090 203360 89140
rect 203140 89020 203150 89090
rect 203350 89020 203360 89090
rect 203140 88980 203360 89020
rect 203140 88910 203150 88980
rect 203350 88910 203360 88980
rect 203140 88860 203360 88910
rect 203640 89090 203860 89140
rect 203640 89020 203650 89090
rect 203850 89020 203860 89090
rect 203640 88980 203860 89020
rect 203640 88910 203650 88980
rect 203850 88910 203860 88980
rect 203640 88860 203860 88910
rect 204140 89090 204360 89140
rect 204140 89020 204150 89090
rect 204350 89020 204360 89090
rect 204140 88980 204360 89020
rect 204140 88910 204150 88980
rect 204350 88910 204360 88980
rect 204140 88860 204360 88910
rect 204640 89090 204860 89140
rect 204640 89020 204650 89090
rect 204850 89020 204860 89090
rect 204640 88980 204860 89020
rect 204640 88910 204650 88980
rect 204850 88910 204860 88980
rect 204640 88860 204860 88910
rect 205140 89090 205360 89140
rect 205140 89020 205150 89090
rect 205350 89020 205360 89090
rect 205140 88980 205360 89020
rect 205140 88910 205150 88980
rect 205350 88910 205360 88980
rect 205140 88860 205360 88910
rect 205640 89090 205860 89140
rect 205640 89020 205650 89090
rect 205850 89020 205860 89090
rect 205640 88980 205860 89020
rect 205640 88910 205650 88980
rect 205850 88910 205860 88980
rect 205640 88860 205860 88910
rect 206140 89090 206360 89140
rect 206140 89020 206150 89090
rect 206350 89020 206360 89090
rect 206140 88980 206360 89020
rect 206140 88910 206150 88980
rect 206350 88910 206360 88980
rect 206140 88860 206360 88910
rect 206640 89090 206860 89140
rect 206640 89020 206650 89090
rect 206850 89020 206860 89090
rect 206640 88980 206860 89020
rect 206640 88910 206650 88980
rect 206850 88910 206860 88980
rect 206640 88860 206860 88910
rect 207140 89090 207360 89140
rect 207140 89020 207150 89090
rect 207350 89020 207360 89090
rect 207140 88980 207360 89020
rect 207140 88910 207150 88980
rect 207350 88910 207360 88980
rect 207140 88860 207360 88910
rect 207640 89090 207860 89140
rect 207640 89020 207650 89090
rect 207850 89020 207860 89090
rect 207640 88980 207860 89020
rect 207640 88910 207650 88980
rect 207850 88910 207860 88980
rect 207640 88860 207860 88910
rect 196000 88850 208000 88860
rect 196000 88650 196020 88850
rect 196090 88650 196410 88850
rect 196480 88650 196520 88850
rect 196590 88650 196910 88850
rect 196980 88650 197020 88850
rect 197090 88650 197410 88850
rect 197480 88650 197520 88850
rect 197590 88650 197910 88850
rect 197980 88650 198020 88850
rect 198090 88650 198410 88850
rect 198480 88650 198520 88850
rect 198590 88650 198910 88850
rect 198980 88650 199020 88850
rect 199090 88650 199410 88850
rect 199480 88650 199520 88850
rect 199590 88650 199910 88850
rect 199980 88650 200020 88850
rect 200090 88650 200410 88850
rect 200480 88650 200520 88850
rect 200590 88650 200910 88850
rect 200980 88650 201020 88850
rect 201090 88650 201410 88850
rect 201480 88650 201520 88850
rect 201590 88650 201910 88850
rect 201980 88650 202020 88850
rect 202090 88650 202410 88850
rect 202480 88650 202520 88850
rect 202590 88650 202910 88850
rect 202980 88650 203020 88850
rect 203090 88650 203410 88850
rect 203480 88650 203520 88850
rect 203590 88650 203910 88850
rect 203980 88650 204020 88850
rect 204090 88650 204410 88850
rect 204480 88650 204520 88850
rect 204590 88650 204910 88850
rect 204980 88650 205020 88850
rect 205090 88650 205410 88850
rect 205480 88650 205520 88850
rect 205590 88650 205910 88850
rect 205980 88650 206020 88850
rect 206090 88650 206410 88850
rect 206480 88650 206520 88850
rect 206590 88650 206910 88850
rect 206980 88650 207020 88850
rect 207090 88650 207410 88850
rect 207480 88650 207520 88850
rect 207590 88650 207910 88850
rect 207980 88650 208000 88850
rect 196000 88640 208000 88650
rect 196140 88590 196360 88640
rect 196140 88520 196150 88590
rect 196350 88520 196360 88590
rect 196140 88480 196360 88520
rect 196140 88410 196150 88480
rect 196350 88410 196360 88480
rect 196140 88360 196360 88410
rect 196640 88590 196860 88640
rect 196640 88520 196650 88590
rect 196850 88520 196860 88590
rect 196640 88480 196860 88520
rect 196640 88410 196650 88480
rect 196850 88410 196860 88480
rect 196640 88360 196860 88410
rect 197140 88590 197360 88640
rect 197140 88520 197150 88590
rect 197350 88520 197360 88590
rect 197140 88480 197360 88520
rect 197140 88410 197150 88480
rect 197350 88410 197360 88480
rect 197140 88360 197360 88410
rect 197640 88590 197860 88640
rect 197640 88520 197650 88590
rect 197850 88520 197860 88590
rect 197640 88480 197860 88520
rect 197640 88410 197650 88480
rect 197850 88410 197860 88480
rect 197640 88360 197860 88410
rect 198140 88590 198360 88640
rect 198140 88520 198150 88590
rect 198350 88520 198360 88590
rect 198140 88480 198360 88520
rect 198140 88410 198150 88480
rect 198350 88410 198360 88480
rect 198140 88360 198360 88410
rect 198640 88590 198860 88640
rect 198640 88520 198650 88590
rect 198850 88520 198860 88590
rect 198640 88480 198860 88520
rect 198640 88410 198650 88480
rect 198850 88410 198860 88480
rect 198640 88360 198860 88410
rect 199140 88590 199360 88640
rect 199140 88520 199150 88590
rect 199350 88520 199360 88590
rect 199140 88480 199360 88520
rect 199140 88410 199150 88480
rect 199350 88410 199360 88480
rect 199140 88360 199360 88410
rect 199640 88590 199860 88640
rect 199640 88520 199650 88590
rect 199850 88520 199860 88590
rect 199640 88480 199860 88520
rect 199640 88410 199650 88480
rect 199850 88410 199860 88480
rect 199640 88360 199860 88410
rect 200140 88590 200360 88640
rect 200140 88520 200150 88590
rect 200350 88520 200360 88590
rect 200140 88480 200360 88520
rect 200140 88410 200150 88480
rect 200350 88410 200360 88480
rect 200140 88360 200360 88410
rect 200640 88590 200860 88640
rect 200640 88520 200650 88590
rect 200850 88520 200860 88590
rect 200640 88480 200860 88520
rect 200640 88410 200650 88480
rect 200850 88410 200860 88480
rect 200640 88360 200860 88410
rect 201140 88590 201360 88640
rect 201140 88520 201150 88590
rect 201350 88520 201360 88590
rect 201140 88480 201360 88520
rect 201140 88410 201150 88480
rect 201350 88410 201360 88480
rect 201140 88360 201360 88410
rect 201640 88590 201860 88640
rect 201640 88520 201650 88590
rect 201850 88520 201860 88590
rect 201640 88480 201860 88520
rect 201640 88410 201650 88480
rect 201850 88410 201860 88480
rect 201640 88360 201860 88410
rect 202140 88590 202360 88640
rect 202140 88520 202150 88590
rect 202350 88520 202360 88590
rect 202140 88480 202360 88520
rect 202140 88410 202150 88480
rect 202350 88410 202360 88480
rect 202140 88360 202360 88410
rect 202640 88590 202860 88640
rect 202640 88520 202650 88590
rect 202850 88520 202860 88590
rect 202640 88480 202860 88520
rect 202640 88410 202650 88480
rect 202850 88410 202860 88480
rect 202640 88360 202860 88410
rect 203140 88590 203360 88640
rect 203140 88520 203150 88590
rect 203350 88520 203360 88590
rect 203140 88480 203360 88520
rect 203140 88410 203150 88480
rect 203350 88410 203360 88480
rect 203140 88360 203360 88410
rect 203640 88590 203860 88640
rect 203640 88520 203650 88590
rect 203850 88520 203860 88590
rect 203640 88480 203860 88520
rect 203640 88410 203650 88480
rect 203850 88410 203860 88480
rect 203640 88360 203860 88410
rect 204140 88590 204360 88640
rect 204140 88520 204150 88590
rect 204350 88520 204360 88590
rect 204140 88480 204360 88520
rect 204140 88410 204150 88480
rect 204350 88410 204360 88480
rect 204140 88360 204360 88410
rect 204640 88590 204860 88640
rect 204640 88520 204650 88590
rect 204850 88520 204860 88590
rect 204640 88480 204860 88520
rect 204640 88410 204650 88480
rect 204850 88410 204860 88480
rect 204640 88360 204860 88410
rect 205140 88590 205360 88640
rect 205140 88520 205150 88590
rect 205350 88520 205360 88590
rect 205140 88480 205360 88520
rect 205140 88410 205150 88480
rect 205350 88410 205360 88480
rect 205140 88360 205360 88410
rect 205640 88590 205860 88640
rect 205640 88520 205650 88590
rect 205850 88520 205860 88590
rect 205640 88480 205860 88520
rect 205640 88410 205650 88480
rect 205850 88410 205860 88480
rect 205640 88360 205860 88410
rect 206140 88590 206360 88640
rect 206140 88520 206150 88590
rect 206350 88520 206360 88590
rect 206140 88480 206360 88520
rect 206140 88410 206150 88480
rect 206350 88410 206360 88480
rect 206140 88360 206360 88410
rect 206640 88590 206860 88640
rect 206640 88520 206650 88590
rect 206850 88520 206860 88590
rect 206640 88480 206860 88520
rect 206640 88410 206650 88480
rect 206850 88410 206860 88480
rect 206640 88360 206860 88410
rect 207140 88590 207360 88640
rect 207140 88520 207150 88590
rect 207350 88520 207360 88590
rect 207140 88480 207360 88520
rect 207140 88410 207150 88480
rect 207350 88410 207360 88480
rect 207140 88360 207360 88410
rect 207640 88590 207860 88640
rect 207640 88520 207650 88590
rect 207850 88520 207860 88590
rect 207640 88480 207860 88520
rect 207640 88410 207650 88480
rect 207850 88410 207860 88480
rect 207640 88360 207860 88410
rect 196000 88350 208000 88360
rect 196000 88150 196020 88350
rect 196090 88150 196410 88350
rect 196480 88150 196520 88350
rect 196590 88150 196910 88350
rect 196980 88150 197020 88350
rect 197090 88150 197410 88350
rect 197480 88150 197520 88350
rect 197590 88150 197910 88350
rect 197980 88150 198020 88350
rect 198090 88150 198410 88350
rect 198480 88150 198520 88350
rect 198590 88150 198910 88350
rect 198980 88150 199020 88350
rect 199090 88150 199410 88350
rect 199480 88150 199520 88350
rect 199590 88150 199910 88350
rect 199980 88150 200020 88350
rect 200090 88150 200410 88350
rect 200480 88150 200520 88350
rect 200590 88150 200910 88350
rect 200980 88150 201020 88350
rect 201090 88150 201410 88350
rect 201480 88150 201520 88350
rect 201590 88150 201910 88350
rect 201980 88150 202020 88350
rect 202090 88150 202410 88350
rect 202480 88150 202520 88350
rect 202590 88150 202910 88350
rect 202980 88150 203020 88350
rect 203090 88150 203410 88350
rect 203480 88150 203520 88350
rect 203590 88150 203910 88350
rect 203980 88150 204020 88350
rect 204090 88150 204410 88350
rect 204480 88150 204520 88350
rect 204590 88150 204910 88350
rect 204980 88150 205020 88350
rect 205090 88150 205410 88350
rect 205480 88150 205520 88350
rect 205590 88150 205910 88350
rect 205980 88150 206020 88350
rect 206090 88150 206410 88350
rect 206480 88150 206520 88350
rect 206590 88150 206910 88350
rect 206980 88150 207020 88350
rect 207090 88150 207410 88350
rect 207480 88150 207520 88350
rect 207590 88150 207910 88350
rect 207980 88150 208000 88350
rect 196000 88140 208000 88150
rect 196140 88090 196360 88140
rect 196140 88020 196150 88090
rect 196350 88020 196360 88090
rect 196140 87980 196360 88020
rect 196140 87910 196150 87980
rect 196350 87910 196360 87980
rect 196140 87860 196360 87910
rect 196640 88090 196860 88140
rect 196640 88020 196650 88090
rect 196850 88020 196860 88090
rect 196640 87980 196860 88020
rect 196640 87910 196650 87980
rect 196850 87910 196860 87980
rect 196640 87860 196860 87910
rect 197140 88090 197360 88140
rect 197140 88020 197150 88090
rect 197350 88020 197360 88090
rect 197140 87980 197360 88020
rect 197140 87910 197150 87980
rect 197350 87910 197360 87980
rect 197140 87860 197360 87910
rect 197640 88090 197860 88140
rect 197640 88020 197650 88090
rect 197850 88020 197860 88090
rect 197640 87980 197860 88020
rect 197640 87910 197650 87980
rect 197850 87910 197860 87980
rect 197640 87860 197860 87910
rect 198140 88090 198360 88140
rect 198140 88020 198150 88090
rect 198350 88020 198360 88090
rect 198140 87980 198360 88020
rect 198140 87910 198150 87980
rect 198350 87910 198360 87980
rect 198140 87860 198360 87910
rect 198640 88090 198860 88140
rect 198640 88020 198650 88090
rect 198850 88020 198860 88090
rect 198640 87980 198860 88020
rect 198640 87910 198650 87980
rect 198850 87910 198860 87980
rect 198640 87860 198860 87910
rect 199140 88090 199360 88140
rect 199140 88020 199150 88090
rect 199350 88020 199360 88090
rect 199140 87980 199360 88020
rect 199140 87910 199150 87980
rect 199350 87910 199360 87980
rect 199140 87860 199360 87910
rect 199640 88090 199860 88140
rect 199640 88020 199650 88090
rect 199850 88020 199860 88090
rect 199640 87980 199860 88020
rect 199640 87910 199650 87980
rect 199850 87910 199860 87980
rect 199640 87860 199860 87910
rect 200140 88090 200360 88140
rect 200140 88020 200150 88090
rect 200350 88020 200360 88090
rect 200140 87980 200360 88020
rect 200140 87910 200150 87980
rect 200350 87910 200360 87980
rect 200140 87860 200360 87910
rect 200640 88090 200860 88140
rect 200640 88020 200650 88090
rect 200850 88020 200860 88090
rect 200640 87980 200860 88020
rect 200640 87910 200650 87980
rect 200850 87910 200860 87980
rect 200640 87860 200860 87910
rect 201140 88090 201360 88140
rect 201140 88020 201150 88090
rect 201350 88020 201360 88090
rect 201140 87980 201360 88020
rect 201140 87910 201150 87980
rect 201350 87910 201360 87980
rect 201140 87860 201360 87910
rect 201640 88090 201860 88140
rect 201640 88020 201650 88090
rect 201850 88020 201860 88090
rect 201640 87980 201860 88020
rect 201640 87910 201650 87980
rect 201850 87910 201860 87980
rect 201640 87860 201860 87910
rect 202140 88090 202360 88140
rect 202140 88020 202150 88090
rect 202350 88020 202360 88090
rect 202140 87980 202360 88020
rect 202140 87910 202150 87980
rect 202350 87910 202360 87980
rect 202140 87860 202360 87910
rect 202640 88090 202860 88140
rect 202640 88020 202650 88090
rect 202850 88020 202860 88090
rect 202640 87980 202860 88020
rect 202640 87910 202650 87980
rect 202850 87910 202860 87980
rect 202640 87860 202860 87910
rect 203140 88090 203360 88140
rect 203140 88020 203150 88090
rect 203350 88020 203360 88090
rect 203140 87980 203360 88020
rect 203140 87910 203150 87980
rect 203350 87910 203360 87980
rect 203140 87860 203360 87910
rect 203640 88090 203860 88140
rect 203640 88020 203650 88090
rect 203850 88020 203860 88090
rect 203640 87980 203860 88020
rect 203640 87910 203650 87980
rect 203850 87910 203860 87980
rect 203640 87860 203860 87910
rect 204140 88090 204360 88140
rect 204140 88020 204150 88090
rect 204350 88020 204360 88090
rect 204140 87980 204360 88020
rect 204140 87910 204150 87980
rect 204350 87910 204360 87980
rect 204140 87860 204360 87910
rect 204640 88090 204860 88140
rect 204640 88020 204650 88090
rect 204850 88020 204860 88090
rect 204640 87980 204860 88020
rect 204640 87910 204650 87980
rect 204850 87910 204860 87980
rect 204640 87860 204860 87910
rect 205140 88090 205360 88140
rect 205140 88020 205150 88090
rect 205350 88020 205360 88090
rect 205140 87980 205360 88020
rect 205140 87910 205150 87980
rect 205350 87910 205360 87980
rect 205140 87860 205360 87910
rect 205640 88090 205860 88140
rect 205640 88020 205650 88090
rect 205850 88020 205860 88090
rect 205640 87980 205860 88020
rect 205640 87910 205650 87980
rect 205850 87910 205860 87980
rect 205640 87860 205860 87910
rect 206140 88090 206360 88140
rect 206140 88020 206150 88090
rect 206350 88020 206360 88090
rect 206140 87980 206360 88020
rect 206140 87910 206150 87980
rect 206350 87910 206360 87980
rect 206140 87860 206360 87910
rect 206640 88090 206860 88140
rect 206640 88020 206650 88090
rect 206850 88020 206860 88090
rect 206640 87980 206860 88020
rect 206640 87910 206650 87980
rect 206850 87910 206860 87980
rect 206640 87860 206860 87910
rect 207140 88090 207360 88140
rect 207140 88020 207150 88090
rect 207350 88020 207360 88090
rect 207140 87980 207360 88020
rect 207140 87910 207150 87980
rect 207350 87910 207360 87980
rect 207140 87860 207360 87910
rect 207640 88090 207860 88140
rect 207640 88020 207650 88090
rect 207850 88020 207860 88090
rect 207640 87980 207860 88020
rect 207640 87910 207650 87980
rect 207850 87910 207860 87980
rect 207640 87860 207860 87910
rect 196000 87850 208000 87860
rect 196000 87650 196020 87850
rect 196090 87650 196410 87850
rect 196480 87650 196520 87850
rect 196590 87650 196910 87850
rect 196980 87650 197020 87850
rect 197090 87650 197410 87850
rect 197480 87650 197520 87850
rect 197590 87650 197910 87850
rect 197980 87650 198020 87850
rect 198090 87650 198410 87850
rect 198480 87650 198520 87850
rect 198590 87650 198910 87850
rect 198980 87650 199020 87850
rect 199090 87650 199410 87850
rect 199480 87650 199520 87850
rect 199590 87650 199910 87850
rect 199980 87650 200020 87850
rect 200090 87650 200410 87850
rect 200480 87650 200520 87850
rect 200590 87650 200910 87850
rect 200980 87650 201020 87850
rect 201090 87650 201410 87850
rect 201480 87650 201520 87850
rect 201590 87650 201910 87850
rect 201980 87650 202020 87850
rect 202090 87650 202410 87850
rect 202480 87650 202520 87850
rect 202590 87650 202910 87850
rect 202980 87650 203020 87850
rect 203090 87650 203410 87850
rect 203480 87650 203520 87850
rect 203590 87650 203910 87850
rect 203980 87650 204020 87850
rect 204090 87650 204410 87850
rect 204480 87650 204520 87850
rect 204590 87650 204910 87850
rect 204980 87650 205020 87850
rect 205090 87650 205410 87850
rect 205480 87650 205520 87850
rect 205590 87650 205910 87850
rect 205980 87650 206020 87850
rect 206090 87650 206410 87850
rect 206480 87650 206520 87850
rect 206590 87650 206910 87850
rect 206980 87650 207020 87850
rect 207090 87650 207410 87850
rect 207480 87650 207520 87850
rect 207590 87650 207910 87850
rect 207980 87650 208000 87850
rect 196000 87640 208000 87650
rect 196140 87590 196360 87640
rect 196140 87520 196150 87590
rect 196350 87520 196360 87590
rect 196140 87480 196360 87520
rect 196140 87410 196150 87480
rect 196350 87410 196360 87480
rect 196140 87360 196360 87410
rect 196640 87590 196860 87640
rect 196640 87520 196650 87590
rect 196850 87520 196860 87590
rect 196640 87480 196860 87520
rect 196640 87410 196650 87480
rect 196850 87410 196860 87480
rect 196640 87360 196860 87410
rect 197140 87590 197360 87640
rect 197140 87520 197150 87590
rect 197350 87520 197360 87590
rect 197140 87480 197360 87520
rect 197140 87410 197150 87480
rect 197350 87410 197360 87480
rect 197140 87360 197360 87410
rect 197640 87590 197860 87640
rect 197640 87520 197650 87590
rect 197850 87520 197860 87590
rect 197640 87480 197860 87520
rect 197640 87410 197650 87480
rect 197850 87410 197860 87480
rect 197640 87360 197860 87410
rect 198140 87590 198360 87640
rect 198140 87520 198150 87590
rect 198350 87520 198360 87590
rect 198140 87480 198360 87520
rect 198140 87410 198150 87480
rect 198350 87410 198360 87480
rect 198140 87360 198360 87410
rect 198640 87590 198860 87640
rect 198640 87520 198650 87590
rect 198850 87520 198860 87590
rect 198640 87480 198860 87520
rect 198640 87410 198650 87480
rect 198850 87410 198860 87480
rect 198640 87360 198860 87410
rect 199140 87590 199360 87640
rect 199140 87520 199150 87590
rect 199350 87520 199360 87590
rect 199140 87480 199360 87520
rect 199140 87410 199150 87480
rect 199350 87410 199360 87480
rect 199140 87360 199360 87410
rect 199640 87590 199860 87640
rect 199640 87520 199650 87590
rect 199850 87520 199860 87590
rect 199640 87480 199860 87520
rect 199640 87410 199650 87480
rect 199850 87410 199860 87480
rect 199640 87360 199860 87410
rect 200140 87590 200360 87640
rect 200140 87520 200150 87590
rect 200350 87520 200360 87590
rect 200140 87480 200360 87520
rect 200140 87410 200150 87480
rect 200350 87410 200360 87480
rect 200140 87360 200360 87410
rect 200640 87590 200860 87640
rect 200640 87520 200650 87590
rect 200850 87520 200860 87590
rect 200640 87480 200860 87520
rect 200640 87410 200650 87480
rect 200850 87410 200860 87480
rect 200640 87360 200860 87410
rect 201140 87590 201360 87640
rect 201140 87520 201150 87590
rect 201350 87520 201360 87590
rect 201140 87480 201360 87520
rect 201140 87410 201150 87480
rect 201350 87410 201360 87480
rect 201140 87360 201360 87410
rect 201640 87590 201860 87640
rect 201640 87520 201650 87590
rect 201850 87520 201860 87590
rect 201640 87480 201860 87520
rect 201640 87410 201650 87480
rect 201850 87410 201860 87480
rect 201640 87360 201860 87410
rect 202140 87590 202360 87640
rect 202140 87520 202150 87590
rect 202350 87520 202360 87590
rect 202140 87480 202360 87520
rect 202140 87410 202150 87480
rect 202350 87410 202360 87480
rect 202140 87360 202360 87410
rect 202640 87590 202860 87640
rect 202640 87520 202650 87590
rect 202850 87520 202860 87590
rect 202640 87480 202860 87520
rect 202640 87410 202650 87480
rect 202850 87410 202860 87480
rect 202640 87360 202860 87410
rect 203140 87590 203360 87640
rect 203140 87520 203150 87590
rect 203350 87520 203360 87590
rect 203140 87480 203360 87520
rect 203140 87410 203150 87480
rect 203350 87410 203360 87480
rect 203140 87360 203360 87410
rect 203640 87590 203860 87640
rect 203640 87520 203650 87590
rect 203850 87520 203860 87590
rect 203640 87480 203860 87520
rect 203640 87410 203650 87480
rect 203850 87410 203860 87480
rect 203640 87360 203860 87410
rect 204140 87590 204360 87640
rect 204140 87520 204150 87590
rect 204350 87520 204360 87590
rect 204140 87480 204360 87520
rect 204140 87410 204150 87480
rect 204350 87410 204360 87480
rect 204140 87360 204360 87410
rect 204640 87590 204860 87640
rect 204640 87520 204650 87590
rect 204850 87520 204860 87590
rect 204640 87480 204860 87520
rect 204640 87410 204650 87480
rect 204850 87410 204860 87480
rect 204640 87360 204860 87410
rect 205140 87590 205360 87640
rect 205140 87520 205150 87590
rect 205350 87520 205360 87590
rect 205140 87480 205360 87520
rect 205140 87410 205150 87480
rect 205350 87410 205360 87480
rect 205140 87360 205360 87410
rect 205640 87590 205860 87640
rect 205640 87520 205650 87590
rect 205850 87520 205860 87590
rect 205640 87480 205860 87520
rect 205640 87410 205650 87480
rect 205850 87410 205860 87480
rect 205640 87360 205860 87410
rect 206140 87590 206360 87640
rect 206140 87520 206150 87590
rect 206350 87520 206360 87590
rect 206140 87480 206360 87520
rect 206140 87410 206150 87480
rect 206350 87410 206360 87480
rect 206140 87360 206360 87410
rect 206640 87590 206860 87640
rect 206640 87520 206650 87590
rect 206850 87520 206860 87590
rect 206640 87480 206860 87520
rect 206640 87410 206650 87480
rect 206850 87410 206860 87480
rect 206640 87360 206860 87410
rect 207140 87590 207360 87640
rect 207140 87520 207150 87590
rect 207350 87520 207360 87590
rect 207140 87480 207360 87520
rect 207140 87410 207150 87480
rect 207350 87410 207360 87480
rect 207140 87360 207360 87410
rect 207640 87590 207860 87640
rect 207640 87520 207650 87590
rect 207850 87520 207860 87590
rect 207640 87480 207860 87520
rect 207640 87410 207650 87480
rect 207850 87410 207860 87480
rect 207640 87360 207860 87410
rect 196000 87350 208000 87360
rect 196000 87150 196020 87350
rect 196090 87150 196410 87350
rect 196480 87150 196520 87350
rect 196590 87150 196910 87350
rect 196980 87150 197020 87350
rect 197090 87150 197410 87350
rect 197480 87150 197520 87350
rect 197590 87150 197910 87350
rect 197980 87150 198020 87350
rect 198090 87150 198410 87350
rect 198480 87150 198520 87350
rect 198590 87150 198910 87350
rect 198980 87150 199020 87350
rect 199090 87150 199410 87350
rect 199480 87150 199520 87350
rect 199590 87150 199910 87350
rect 199980 87150 200020 87350
rect 200090 87150 200410 87350
rect 200480 87150 200520 87350
rect 200590 87150 200910 87350
rect 200980 87150 201020 87350
rect 201090 87150 201410 87350
rect 201480 87150 201520 87350
rect 201590 87150 201910 87350
rect 201980 87150 202020 87350
rect 202090 87150 202410 87350
rect 202480 87150 202520 87350
rect 202590 87150 202910 87350
rect 202980 87150 203020 87350
rect 203090 87150 203410 87350
rect 203480 87150 203520 87350
rect 203590 87150 203910 87350
rect 203980 87150 204020 87350
rect 204090 87150 204410 87350
rect 204480 87150 204520 87350
rect 204590 87150 204910 87350
rect 204980 87150 205020 87350
rect 205090 87150 205410 87350
rect 205480 87150 205520 87350
rect 205590 87150 205910 87350
rect 205980 87150 206020 87350
rect 206090 87150 206410 87350
rect 206480 87150 206520 87350
rect 206590 87150 206910 87350
rect 206980 87150 207020 87350
rect 207090 87150 207410 87350
rect 207480 87150 207520 87350
rect 207590 87150 207910 87350
rect 207980 87150 208000 87350
rect 196000 87140 208000 87150
rect 128750 87110 128910 87120
rect 128750 86870 128760 87110
rect 128900 86870 128910 87110
rect 128750 86860 128910 86870
rect 129070 87110 129230 87120
rect 129070 86870 129080 87110
rect 129220 86870 129230 87110
rect 129070 86860 129230 86870
rect 196140 87090 196360 87140
rect 196140 87020 196150 87090
rect 196350 87020 196360 87090
rect 196140 86980 196360 87020
rect 196140 86910 196150 86980
rect 196350 86910 196360 86980
rect 196140 86860 196360 86910
rect 196640 87090 196860 87140
rect 196640 87020 196650 87090
rect 196850 87020 196860 87090
rect 196640 86980 196860 87020
rect 196640 86910 196650 86980
rect 196850 86910 196860 86980
rect 196640 86860 196860 86910
rect 197140 87090 197360 87140
rect 197140 87020 197150 87090
rect 197350 87020 197360 87090
rect 197140 86980 197360 87020
rect 197140 86910 197150 86980
rect 197350 86910 197360 86980
rect 197140 86860 197360 86910
rect 197640 87090 197860 87140
rect 197640 87020 197650 87090
rect 197850 87020 197860 87090
rect 197640 86980 197860 87020
rect 197640 86910 197650 86980
rect 197850 86910 197860 86980
rect 197640 86860 197860 86910
rect 198140 87090 198360 87140
rect 198140 87020 198150 87090
rect 198350 87020 198360 87090
rect 198140 86980 198360 87020
rect 198140 86910 198150 86980
rect 198350 86910 198360 86980
rect 198140 86860 198360 86910
rect 198640 87090 198860 87140
rect 198640 87020 198650 87090
rect 198850 87020 198860 87090
rect 198640 86980 198860 87020
rect 198640 86910 198650 86980
rect 198850 86910 198860 86980
rect 198640 86860 198860 86910
rect 199140 87090 199360 87140
rect 199140 87020 199150 87090
rect 199350 87020 199360 87090
rect 199140 86980 199360 87020
rect 199140 86910 199150 86980
rect 199350 86910 199360 86980
rect 199140 86860 199360 86910
rect 199640 87090 199860 87140
rect 199640 87020 199650 87090
rect 199850 87020 199860 87090
rect 199640 86980 199860 87020
rect 199640 86910 199650 86980
rect 199850 86910 199860 86980
rect 199640 86860 199860 86910
rect 200140 87090 200360 87140
rect 200140 87020 200150 87090
rect 200350 87020 200360 87090
rect 200140 86980 200360 87020
rect 200140 86910 200150 86980
rect 200350 86910 200360 86980
rect 200140 86860 200360 86910
rect 200640 87090 200860 87140
rect 200640 87020 200650 87090
rect 200850 87020 200860 87090
rect 200640 86980 200860 87020
rect 200640 86910 200650 86980
rect 200850 86910 200860 86980
rect 200640 86860 200860 86910
rect 201140 87090 201360 87140
rect 201140 87020 201150 87090
rect 201350 87020 201360 87090
rect 201140 86980 201360 87020
rect 201140 86910 201150 86980
rect 201350 86910 201360 86980
rect 201140 86860 201360 86910
rect 201640 87090 201860 87140
rect 201640 87020 201650 87090
rect 201850 87020 201860 87090
rect 201640 86980 201860 87020
rect 201640 86910 201650 86980
rect 201850 86910 201860 86980
rect 201640 86860 201860 86910
rect 202140 87090 202360 87140
rect 202140 87020 202150 87090
rect 202350 87020 202360 87090
rect 202140 86980 202360 87020
rect 202140 86910 202150 86980
rect 202350 86910 202360 86980
rect 202140 86860 202360 86910
rect 202640 87090 202860 87140
rect 202640 87020 202650 87090
rect 202850 87020 202860 87090
rect 202640 86980 202860 87020
rect 202640 86910 202650 86980
rect 202850 86910 202860 86980
rect 202640 86860 202860 86910
rect 203140 87090 203360 87140
rect 203140 87020 203150 87090
rect 203350 87020 203360 87090
rect 203140 86980 203360 87020
rect 203140 86910 203150 86980
rect 203350 86910 203360 86980
rect 203140 86860 203360 86910
rect 203640 87090 203860 87140
rect 203640 87020 203650 87090
rect 203850 87020 203860 87090
rect 203640 86980 203860 87020
rect 203640 86910 203650 86980
rect 203850 86910 203860 86980
rect 203640 86860 203860 86910
rect 204140 87090 204360 87140
rect 204140 87020 204150 87090
rect 204350 87020 204360 87090
rect 204140 86980 204360 87020
rect 204140 86910 204150 86980
rect 204350 86910 204360 86980
rect 204140 86860 204360 86910
rect 204640 87090 204860 87140
rect 204640 87020 204650 87090
rect 204850 87020 204860 87090
rect 204640 86980 204860 87020
rect 204640 86910 204650 86980
rect 204850 86910 204860 86980
rect 204640 86860 204860 86910
rect 205140 87090 205360 87140
rect 205140 87020 205150 87090
rect 205350 87020 205360 87090
rect 205140 86980 205360 87020
rect 205140 86910 205150 86980
rect 205350 86910 205360 86980
rect 205140 86860 205360 86910
rect 205640 87090 205860 87140
rect 205640 87020 205650 87090
rect 205850 87020 205860 87090
rect 205640 86980 205860 87020
rect 205640 86910 205650 86980
rect 205850 86910 205860 86980
rect 205640 86860 205860 86910
rect 206140 87090 206360 87140
rect 206140 87020 206150 87090
rect 206350 87020 206360 87090
rect 206140 86980 206360 87020
rect 206140 86910 206150 86980
rect 206350 86910 206360 86980
rect 206140 86860 206360 86910
rect 206640 87090 206860 87140
rect 206640 87020 206650 87090
rect 206850 87020 206860 87090
rect 206640 86980 206860 87020
rect 206640 86910 206650 86980
rect 206850 86910 206860 86980
rect 206640 86860 206860 86910
rect 207140 87090 207360 87140
rect 207140 87020 207150 87090
rect 207350 87020 207360 87090
rect 207140 86980 207360 87020
rect 207140 86910 207150 86980
rect 207350 86910 207360 86980
rect 207140 86860 207360 86910
rect 207640 87090 207860 87140
rect 207640 87020 207650 87090
rect 207850 87020 207860 87090
rect 207640 86980 207860 87020
rect 207640 86910 207650 86980
rect 207850 86910 207860 86980
rect 207640 86860 207860 86910
rect 196000 86850 208000 86860
rect 196000 86650 196020 86850
rect 196090 86650 196410 86850
rect 196480 86650 196520 86850
rect 196590 86650 196910 86850
rect 196980 86650 197020 86850
rect 197090 86650 197410 86850
rect 197480 86650 197520 86850
rect 197590 86650 197910 86850
rect 197980 86650 198020 86850
rect 198090 86650 198410 86850
rect 198480 86650 198520 86850
rect 198590 86650 198910 86850
rect 198980 86650 199020 86850
rect 199090 86650 199410 86850
rect 199480 86650 199520 86850
rect 199590 86650 199910 86850
rect 199980 86650 200020 86850
rect 200090 86650 200410 86850
rect 200480 86650 200520 86850
rect 200590 86650 200910 86850
rect 200980 86650 201020 86850
rect 201090 86650 201410 86850
rect 201480 86650 201520 86850
rect 201590 86650 201910 86850
rect 201980 86650 202020 86850
rect 202090 86650 202410 86850
rect 202480 86650 202520 86850
rect 202590 86650 202910 86850
rect 202980 86650 203020 86850
rect 203090 86650 203410 86850
rect 203480 86650 203520 86850
rect 203590 86650 203910 86850
rect 203980 86650 204020 86850
rect 204090 86650 204410 86850
rect 204480 86650 204520 86850
rect 204590 86650 204910 86850
rect 204980 86650 205020 86850
rect 205090 86650 205410 86850
rect 205480 86650 205520 86850
rect 205590 86650 205910 86850
rect 205980 86650 206020 86850
rect 206090 86650 206410 86850
rect 206480 86650 206520 86850
rect 206590 86650 206910 86850
rect 206980 86650 207020 86850
rect 207090 86650 207410 86850
rect 207480 86650 207520 86850
rect 207590 86650 207910 86850
rect 207980 86650 208000 86850
rect 196000 86640 208000 86650
rect 128860 86630 129040 86640
rect 128860 86510 128870 86630
rect 129030 86510 129040 86630
rect 128860 86500 129040 86510
rect 196140 86590 196360 86640
rect 196140 86520 196150 86590
rect 196350 86520 196360 86590
rect 196140 86480 196360 86520
rect 196140 86410 196150 86480
rect 196350 86410 196360 86480
rect 196140 86360 196360 86410
rect 196640 86590 196860 86640
rect 196640 86520 196650 86590
rect 196850 86520 196860 86590
rect 196640 86480 196860 86520
rect 196640 86410 196650 86480
rect 196850 86410 196860 86480
rect 196640 86360 196860 86410
rect 197140 86590 197360 86640
rect 197140 86520 197150 86590
rect 197350 86520 197360 86590
rect 197140 86480 197360 86520
rect 197140 86410 197150 86480
rect 197350 86410 197360 86480
rect 197140 86360 197360 86410
rect 197640 86590 197860 86640
rect 197640 86520 197650 86590
rect 197850 86520 197860 86590
rect 197640 86480 197860 86520
rect 197640 86410 197650 86480
rect 197850 86410 197860 86480
rect 197640 86360 197860 86410
rect 198140 86590 198360 86640
rect 198140 86520 198150 86590
rect 198350 86520 198360 86590
rect 198140 86480 198360 86520
rect 198140 86410 198150 86480
rect 198350 86410 198360 86480
rect 198140 86360 198360 86410
rect 198640 86590 198860 86640
rect 198640 86520 198650 86590
rect 198850 86520 198860 86590
rect 198640 86480 198860 86520
rect 198640 86410 198650 86480
rect 198850 86410 198860 86480
rect 198640 86360 198860 86410
rect 199140 86590 199360 86640
rect 199140 86520 199150 86590
rect 199350 86520 199360 86590
rect 199140 86480 199360 86520
rect 199140 86410 199150 86480
rect 199350 86410 199360 86480
rect 199140 86360 199360 86410
rect 199640 86590 199860 86640
rect 199640 86520 199650 86590
rect 199850 86520 199860 86590
rect 199640 86480 199860 86520
rect 199640 86410 199650 86480
rect 199850 86410 199860 86480
rect 199640 86360 199860 86410
rect 200140 86590 200360 86640
rect 200140 86520 200150 86590
rect 200350 86520 200360 86590
rect 200140 86480 200360 86520
rect 200140 86410 200150 86480
rect 200350 86410 200360 86480
rect 200140 86360 200360 86410
rect 200640 86590 200860 86640
rect 200640 86520 200650 86590
rect 200850 86520 200860 86590
rect 200640 86480 200860 86520
rect 200640 86410 200650 86480
rect 200850 86410 200860 86480
rect 200640 86360 200860 86410
rect 201140 86590 201360 86640
rect 201140 86520 201150 86590
rect 201350 86520 201360 86590
rect 201140 86480 201360 86520
rect 201140 86410 201150 86480
rect 201350 86410 201360 86480
rect 201140 86360 201360 86410
rect 201640 86590 201860 86640
rect 201640 86520 201650 86590
rect 201850 86520 201860 86590
rect 201640 86480 201860 86520
rect 201640 86410 201650 86480
rect 201850 86410 201860 86480
rect 201640 86360 201860 86410
rect 202140 86590 202360 86640
rect 202140 86520 202150 86590
rect 202350 86520 202360 86590
rect 202140 86480 202360 86520
rect 202140 86410 202150 86480
rect 202350 86410 202360 86480
rect 202140 86360 202360 86410
rect 202640 86590 202860 86640
rect 202640 86520 202650 86590
rect 202850 86520 202860 86590
rect 202640 86480 202860 86520
rect 202640 86410 202650 86480
rect 202850 86410 202860 86480
rect 202640 86360 202860 86410
rect 203140 86590 203360 86640
rect 203140 86520 203150 86590
rect 203350 86520 203360 86590
rect 203140 86480 203360 86520
rect 203140 86410 203150 86480
rect 203350 86410 203360 86480
rect 203140 86360 203360 86410
rect 203640 86590 203860 86640
rect 203640 86520 203650 86590
rect 203850 86520 203860 86590
rect 203640 86480 203860 86520
rect 203640 86410 203650 86480
rect 203850 86410 203860 86480
rect 203640 86360 203860 86410
rect 204140 86590 204360 86640
rect 204140 86520 204150 86590
rect 204350 86520 204360 86590
rect 204140 86480 204360 86520
rect 204140 86410 204150 86480
rect 204350 86410 204360 86480
rect 204140 86360 204360 86410
rect 204640 86590 204860 86640
rect 204640 86520 204650 86590
rect 204850 86520 204860 86590
rect 204640 86480 204860 86520
rect 204640 86410 204650 86480
rect 204850 86410 204860 86480
rect 204640 86360 204860 86410
rect 205140 86590 205360 86640
rect 205140 86520 205150 86590
rect 205350 86520 205360 86590
rect 205140 86480 205360 86520
rect 205140 86410 205150 86480
rect 205350 86410 205360 86480
rect 205140 86360 205360 86410
rect 205640 86590 205860 86640
rect 205640 86520 205650 86590
rect 205850 86520 205860 86590
rect 205640 86480 205860 86520
rect 205640 86410 205650 86480
rect 205850 86410 205860 86480
rect 205640 86360 205860 86410
rect 206140 86590 206360 86640
rect 206140 86520 206150 86590
rect 206350 86520 206360 86590
rect 206140 86480 206360 86520
rect 206140 86410 206150 86480
rect 206350 86410 206360 86480
rect 206140 86360 206360 86410
rect 206640 86590 206860 86640
rect 206640 86520 206650 86590
rect 206850 86520 206860 86590
rect 206640 86480 206860 86520
rect 206640 86410 206650 86480
rect 206850 86410 206860 86480
rect 206640 86360 206860 86410
rect 207140 86590 207360 86640
rect 207140 86520 207150 86590
rect 207350 86520 207360 86590
rect 207140 86480 207360 86520
rect 207140 86410 207150 86480
rect 207350 86410 207360 86480
rect 207140 86360 207360 86410
rect 207640 86590 207860 86640
rect 207640 86520 207650 86590
rect 207850 86520 207860 86590
rect 207640 86480 207860 86520
rect 207640 86410 207650 86480
rect 207850 86410 207860 86480
rect 207640 86360 207860 86410
rect 196000 86350 208000 86360
rect 196000 86150 196020 86350
rect 196090 86150 196410 86350
rect 196480 86150 196520 86350
rect 196590 86150 196910 86350
rect 196980 86150 197020 86350
rect 197090 86150 197410 86350
rect 197480 86150 197520 86350
rect 197590 86150 197910 86350
rect 197980 86150 198020 86350
rect 198090 86150 198410 86350
rect 198480 86150 198520 86350
rect 198590 86150 198910 86350
rect 198980 86150 199020 86350
rect 199090 86150 199410 86350
rect 199480 86150 199520 86350
rect 199590 86150 199910 86350
rect 199980 86150 200020 86350
rect 200090 86150 200410 86350
rect 200480 86150 200520 86350
rect 200590 86150 200910 86350
rect 200980 86150 201020 86350
rect 201090 86150 201410 86350
rect 201480 86150 201520 86350
rect 201590 86150 201910 86350
rect 201980 86150 202020 86350
rect 202090 86150 202410 86350
rect 202480 86150 202520 86350
rect 202590 86150 202910 86350
rect 202980 86150 203020 86350
rect 203090 86150 203410 86350
rect 203480 86150 203520 86350
rect 203590 86150 203910 86350
rect 203980 86150 204020 86350
rect 204090 86150 204410 86350
rect 204480 86150 204520 86350
rect 204590 86150 204910 86350
rect 204980 86150 205020 86350
rect 205090 86150 205410 86350
rect 205480 86150 205520 86350
rect 205590 86150 205910 86350
rect 205980 86150 206020 86350
rect 206090 86150 206410 86350
rect 206480 86150 206520 86350
rect 206590 86150 206910 86350
rect 206980 86150 207020 86350
rect 207090 86150 207410 86350
rect 207480 86150 207520 86350
rect 207590 86150 207910 86350
rect 207980 86150 208000 86350
rect 196000 86140 208000 86150
rect 196140 86090 196360 86140
rect 196140 86020 196150 86090
rect 196350 86020 196360 86090
rect 196140 85980 196360 86020
rect 196140 85910 196150 85980
rect 196350 85910 196360 85980
rect 196140 85860 196360 85910
rect 196640 86090 196860 86140
rect 196640 86020 196650 86090
rect 196850 86020 196860 86090
rect 196640 85980 196860 86020
rect 196640 85910 196650 85980
rect 196850 85910 196860 85980
rect 196640 85860 196860 85910
rect 197140 86090 197360 86140
rect 197140 86020 197150 86090
rect 197350 86020 197360 86090
rect 197140 85980 197360 86020
rect 197140 85910 197150 85980
rect 197350 85910 197360 85980
rect 197140 85860 197360 85910
rect 197640 86090 197860 86140
rect 197640 86020 197650 86090
rect 197850 86020 197860 86090
rect 197640 85980 197860 86020
rect 197640 85910 197650 85980
rect 197850 85910 197860 85980
rect 197640 85860 197860 85910
rect 198140 86090 198360 86140
rect 198140 86020 198150 86090
rect 198350 86020 198360 86090
rect 198140 85980 198360 86020
rect 198140 85910 198150 85980
rect 198350 85910 198360 85980
rect 198140 85860 198360 85910
rect 198640 86090 198860 86140
rect 198640 86020 198650 86090
rect 198850 86020 198860 86090
rect 198640 85980 198860 86020
rect 198640 85910 198650 85980
rect 198850 85910 198860 85980
rect 198640 85860 198860 85910
rect 199140 86090 199360 86140
rect 199140 86020 199150 86090
rect 199350 86020 199360 86090
rect 199140 85980 199360 86020
rect 199140 85910 199150 85980
rect 199350 85910 199360 85980
rect 199140 85860 199360 85910
rect 199640 86090 199860 86140
rect 199640 86020 199650 86090
rect 199850 86020 199860 86090
rect 199640 85980 199860 86020
rect 199640 85910 199650 85980
rect 199850 85910 199860 85980
rect 199640 85860 199860 85910
rect 200140 86090 200360 86140
rect 200140 86020 200150 86090
rect 200350 86020 200360 86090
rect 200140 85980 200360 86020
rect 200140 85910 200150 85980
rect 200350 85910 200360 85980
rect 200140 85860 200360 85910
rect 200640 86090 200860 86140
rect 200640 86020 200650 86090
rect 200850 86020 200860 86090
rect 200640 85980 200860 86020
rect 200640 85910 200650 85980
rect 200850 85910 200860 85980
rect 200640 85860 200860 85910
rect 201140 86090 201360 86140
rect 201140 86020 201150 86090
rect 201350 86020 201360 86090
rect 201140 85980 201360 86020
rect 201140 85910 201150 85980
rect 201350 85910 201360 85980
rect 201140 85860 201360 85910
rect 201640 86090 201860 86140
rect 201640 86020 201650 86090
rect 201850 86020 201860 86090
rect 201640 85980 201860 86020
rect 201640 85910 201650 85980
rect 201850 85910 201860 85980
rect 201640 85860 201860 85910
rect 202140 86090 202360 86140
rect 202140 86020 202150 86090
rect 202350 86020 202360 86090
rect 202140 85980 202360 86020
rect 202140 85910 202150 85980
rect 202350 85910 202360 85980
rect 202140 85860 202360 85910
rect 202640 86090 202860 86140
rect 202640 86020 202650 86090
rect 202850 86020 202860 86090
rect 202640 85980 202860 86020
rect 202640 85910 202650 85980
rect 202850 85910 202860 85980
rect 202640 85860 202860 85910
rect 203140 86090 203360 86140
rect 203140 86020 203150 86090
rect 203350 86020 203360 86090
rect 203140 85980 203360 86020
rect 203140 85910 203150 85980
rect 203350 85910 203360 85980
rect 203140 85860 203360 85910
rect 203640 86090 203860 86140
rect 203640 86020 203650 86090
rect 203850 86020 203860 86090
rect 203640 85980 203860 86020
rect 203640 85910 203650 85980
rect 203850 85910 203860 85980
rect 203640 85860 203860 85910
rect 204140 86090 204360 86140
rect 204140 86020 204150 86090
rect 204350 86020 204360 86090
rect 204140 85980 204360 86020
rect 204140 85910 204150 85980
rect 204350 85910 204360 85980
rect 204140 85860 204360 85910
rect 204640 86090 204860 86140
rect 204640 86020 204650 86090
rect 204850 86020 204860 86090
rect 204640 85980 204860 86020
rect 204640 85910 204650 85980
rect 204850 85910 204860 85980
rect 204640 85860 204860 85910
rect 205140 86090 205360 86140
rect 205140 86020 205150 86090
rect 205350 86020 205360 86090
rect 205140 85980 205360 86020
rect 205140 85910 205150 85980
rect 205350 85910 205360 85980
rect 205140 85860 205360 85910
rect 205640 86090 205860 86140
rect 205640 86020 205650 86090
rect 205850 86020 205860 86090
rect 205640 85980 205860 86020
rect 205640 85910 205650 85980
rect 205850 85910 205860 85980
rect 205640 85860 205860 85910
rect 206140 86090 206360 86140
rect 206140 86020 206150 86090
rect 206350 86020 206360 86090
rect 206140 85980 206360 86020
rect 206140 85910 206150 85980
rect 206350 85910 206360 85980
rect 206140 85860 206360 85910
rect 206640 86090 206860 86140
rect 206640 86020 206650 86090
rect 206850 86020 206860 86090
rect 206640 85980 206860 86020
rect 206640 85910 206650 85980
rect 206850 85910 206860 85980
rect 206640 85860 206860 85910
rect 207140 86090 207360 86140
rect 207140 86020 207150 86090
rect 207350 86020 207360 86090
rect 207140 85980 207360 86020
rect 207140 85910 207150 85980
rect 207350 85910 207360 85980
rect 207140 85860 207360 85910
rect 207640 86090 207860 86140
rect 207640 86020 207650 86090
rect 207850 86020 207860 86090
rect 207640 85980 207860 86020
rect 207640 85910 207650 85980
rect 207850 85910 207860 85980
rect 207640 85860 207860 85910
rect 196000 85850 208000 85860
rect 196000 85650 196020 85850
rect 196090 85650 196410 85850
rect 196480 85650 196520 85850
rect 196590 85650 196910 85850
rect 196980 85650 197020 85850
rect 197090 85650 197410 85850
rect 197480 85650 197520 85850
rect 197590 85650 197910 85850
rect 197980 85650 198020 85850
rect 198090 85650 198410 85850
rect 198480 85650 198520 85850
rect 198590 85650 198910 85850
rect 198980 85650 199020 85850
rect 199090 85650 199410 85850
rect 199480 85650 199520 85850
rect 199590 85650 199910 85850
rect 199980 85650 200020 85850
rect 200090 85650 200410 85850
rect 200480 85650 200520 85850
rect 200590 85650 200910 85850
rect 200980 85650 201020 85850
rect 201090 85650 201410 85850
rect 201480 85650 201520 85850
rect 201590 85650 201910 85850
rect 201980 85650 202020 85850
rect 202090 85650 202410 85850
rect 202480 85650 202520 85850
rect 202590 85650 202910 85850
rect 202980 85650 203020 85850
rect 203090 85650 203410 85850
rect 203480 85650 203520 85850
rect 203590 85650 203910 85850
rect 203980 85650 204020 85850
rect 204090 85650 204410 85850
rect 204480 85650 204520 85850
rect 204590 85650 204910 85850
rect 204980 85650 205020 85850
rect 205090 85650 205410 85850
rect 205480 85650 205520 85850
rect 205590 85650 205910 85850
rect 205980 85650 206020 85850
rect 206090 85650 206410 85850
rect 206480 85650 206520 85850
rect 206590 85650 206910 85850
rect 206980 85650 207020 85850
rect 207090 85650 207410 85850
rect 207480 85650 207520 85850
rect 207590 85650 207910 85850
rect 207980 85650 208000 85850
rect 196000 85640 208000 85650
rect 196140 85590 196360 85640
rect 196140 85520 196150 85590
rect 196350 85520 196360 85590
rect 196140 85480 196360 85520
rect 196140 85410 196150 85480
rect 196350 85410 196360 85480
rect 196140 85360 196360 85410
rect 196640 85590 196860 85640
rect 196640 85520 196650 85590
rect 196850 85520 196860 85590
rect 196640 85480 196860 85520
rect 196640 85410 196650 85480
rect 196850 85410 196860 85480
rect 196640 85360 196860 85410
rect 197140 85590 197360 85640
rect 197140 85520 197150 85590
rect 197350 85520 197360 85590
rect 197140 85480 197360 85520
rect 197140 85410 197150 85480
rect 197350 85410 197360 85480
rect 197140 85360 197360 85410
rect 197640 85590 197860 85640
rect 197640 85520 197650 85590
rect 197850 85520 197860 85590
rect 197640 85480 197860 85520
rect 197640 85410 197650 85480
rect 197850 85410 197860 85480
rect 197640 85360 197860 85410
rect 198140 85590 198360 85640
rect 198140 85520 198150 85590
rect 198350 85520 198360 85590
rect 198140 85480 198360 85520
rect 198140 85410 198150 85480
rect 198350 85410 198360 85480
rect 198140 85360 198360 85410
rect 198640 85590 198860 85640
rect 198640 85520 198650 85590
rect 198850 85520 198860 85590
rect 198640 85480 198860 85520
rect 198640 85410 198650 85480
rect 198850 85410 198860 85480
rect 198640 85360 198860 85410
rect 199140 85590 199360 85640
rect 199140 85520 199150 85590
rect 199350 85520 199360 85590
rect 199140 85480 199360 85520
rect 199140 85410 199150 85480
rect 199350 85410 199360 85480
rect 199140 85360 199360 85410
rect 199640 85590 199860 85640
rect 199640 85520 199650 85590
rect 199850 85520 199860 85590
rect 199640 85480 199860 85520
rect 199640 85410 199650 85480
rect 199850 85410 199860 85480
rect 199640 85360 199860 85410
rect 200140 85590 200360 85640
rect 200140 85520 200150 85590
rect 200350 85520 200360 85590
rect 200140 85480 200360 85520
rect 200140 85410 200150 85480
rect 200350 85410 200360 85480
rect 200140 85360 200360 85410
rect 200640 85590 200860 85640
rect 200640 85520 200650 85590
rect 200850 85520 200860 85590
rect 200640 85480 200860 85520
rect 200640 85410 200650 85480
rect 200850 85410 200860 85480
rect 200640 85360 200860 85410
rect 201140 85590 201360 85640
rect 201140 85520 201150 85590
rect 201350 85520 201360 85590
rect 201140 85480 201360 85520
rect 201140 85410 201150 85480
rect 201350 85410 201360 85480
rect 201140 85360 201360 85410
rect 201640 85590 201860 85640
rect 201640 85520 201650 85590
rect 201850 85520 201860 85590
rect 201640 85480 201860 85520
rect 201640 85410 201650 85480
rect 201850 85410 201860 85480
rect 201640 85360 201860 85410
rect 202140 85590 202360 85640
rect 202140 85520 202150 85590
rect 202350 85520 202360 85590
rect 202140 85480 202360 85520
rect 202140 85410 202150 85480
rect 202350 85410 202360 85480
rect 202140 85360 202360 85410
rect 202640 85590 202860 85640
rect 202640 85520 202650 85590
rect 202850 85520 202860 85590
rect 202640 85480 202860 85520
rect 202640 85410 202650 85480
rect 202850 85410 202860 85480
rect 202640 85360 202860 85410
rect 203140 85590 203360 85640
rect 203140 85520 203150 85590
rect 203350 85520 203360 85590
rect 203140 85480 203360 85520
rect 203140 85410 203150 85480
rect 203350 85410 203360 85480
rect 203140 85360 203360 85410
rect 203640 85590 203860 85640
rect 203640 85520 203650 85590
rect 203850 85520 203860 85590
rect 203640 85480 203860 85520
rect 203640 85410 203650 85480
rect 203850 85410 203860 85480
rect 203640 85360 203860 85410
rect 204140 85590 204360 85640
rect 204140 85520 204150 85590
rect 204350 85520 204360 85590
rect 204140 85480 204360 85520
rect 204140 85410 204150 85480
rect 204350 85410 204360 85480
rect 204140 85360 204360 85410
rect 204640 85590 204860 85640
rect 204640 85520 204650 85590
rect 204850 85520 204860 85590
rect 204640 85480 204860 85520
rect 204640 85410 204650 85480
rect 204850 85410 204860 85480
rect 204640 85360 204860 85410
rect 205140 85590 205360 85640
rect 205140 85520 205150 85590
rect 205350 85520 205360 85590
rect 205140 85480 205360 85520
rect 205140 85410 205150 85480
rect 205350 85410 205360 85480
rect 205140 85360 205360 85410
rect 205640 85590 205860 85640
rect 205640 85520 205650 85590
rect 205850 85520 205860 85590
rect 205640 85480 205860 85520
rect 205640 85410 205650 85480
rect 205850 85410 205860 85480
rect 205640 85360 205860 85410
rect 206140 85590 206360 85640
rect 206140 85520 206150 85590
rect 206350 85520 206360 85590
rect 206140 85480 206360 85520
rect 206140 85410 206150 85480
rect 206350 85410 206360 85480
rect 206140 85360 206360 85410
rect 206640 85590 206860 85640
rect 206640 85520 206650 85590
rect 206850 85520 206860 85590
rect 206640 85480 206860 85520
rect 206640 85410 206650 85480
rect 206850 85410 206860 85480
rect 206640 85360 206860 85410
rect 207140 85590 207360 85640
rect 207140 85520 207150 85590
rect 207350 85520 207360 85590
rect 207140 85480 207360 85520
rect 207140 85410 207150 85480
rect 207350 85410 207360 85480
rect 207140 85360 207360 85410
rect 207640 85590 207860 85640
rect 207640 85520 207650 85590
rect 207850 85520 207860 85590
rect 207640 85480 207860 85520
rect 207640 85410 207650 85480
rect 207850 85410 207860 85480
rect 207640 85360 207860 85410
rect 196000 85350 208000 85360
rect 196000 85150 196020 85350
rect 196090 85150 196410 85350
rect 196480 85150 196520 85350
rect 196590 85150 196910 85350
rect 196980 85150 197020 85350
rect 197090 85150 197410 85350
rect 197480 85150 197520 85350
rect 197590 85150 197910 85350
rect 197980 85150 198020 85350
rect 198090 85150 198410 85350
rect 198480 85150 198520 85350
rect 198590 85150 198910 85350
rect 198980 85150 199020 85350
rect 199090 85150 199410 85350
rect 199480 85150 199520 85350
rect 199590 85150 199910 85350
rect 199980 85150 200020 85350
rect 200090 85150 200410 85350
rect 200480 85150 200520 85350
rect 200590 85150 200910 85350
rect 200980 85150 201020 85350
rect 201090 85150 201410 85350
rect 201480 85150 201520 85350
rect 201590 85150 201910 85350
rect 201980 85150 202020 85350
rect 202090 85150 202410 85350
rect 202480 85150 202520 85350
rect 202590 85150 202910 85350
rect 202980 85150 203020 85350
rect 203090 85150 203410 85350
rect 203480 85150 203520 85350
rect 203590 85150 203910 85350
rect 203980 85150 204020 85350
rect 204090 85150 204410 85350
rect 204480 85150 204520 85350
rect 204590 85150 204910 85350
rect 204980 85150 205020 85350
rect 205090 85150 205410 85350
rect 205480 85150 205520 85350
rect 205590 85150 205910 85350
rect 205980 85150 206020 85350
rect 206090 85150 206410 85350
rect 206480 85150 206520 85350
rect 206590 85150 206910 85350
rect 206980 85150 207020 85350
rect 207090 85150 207410 85350
rect 207480 85150 207520 85350
rect 207590 85150 207910 85350
rect 207980 85150 208000 85350
rect 196000 85140 208000 85150
rect 196140 85090 196360 85140
rect 196140 85020 196150 85090
rect 196350 85020 196360 85090
rect 196140 84980 196360 85020
rect 196140 84910 196150 84980
rect 196350 84910 196360 84980
rect 196140 84860 196360 84910
rect 196640 85090 196860 85140
rect 196640 85020 196650 85090
rect 196850 85020 196860 85090
rect 196640 84980 196860 85020
rect 196640 84910 196650 84980
rect 196850 84910 196860 84980
rect 196640 84860 196860 84910
rect 197140 85090 197360 85140
rect 197140 85020 197150 85090
rect 197350 85020 197360 85090
rect 197140 84980 197360 85020
rect 197140 84910 197150 84980
rect 197350 84910 197360 84980
rect 197140 84860 197360 84910
rect 197640 85090 197860 85140
rect 197640 85020 197650 85090
rect 197850 85020 197860 85090
rect 197640 84980 197860 85020
rect 197640 84910 197650 84980
rect 197850 84910 197860 84980
rect 197640 84860 197860 84910
rect 198140 85090 198360 85140
rect 198140 85020 198150 85090
rect 198350 85020 198360 85090
rect 198140 84980 198360 85020
rect 198140 84910 198150 84980
rect 198350 84910 198360 84980
rect 198140 84860 198360 84910
rect 198640 85090 198860 85140
rect 198640 85020 198650 85090
rect 198850 85020 198860 85090
rect 198640 84980 198860 85020
rect 198640 84910 198650 84980
rect 198850 84910 198860 84980
rect 198640 84860 198860 84910
rect 199140 85090 199360 85140
rect 199140 85020 199150 85090
rect 199350 85020 199360 85090
rect 199140 84980 199360 85020
rect 199140 84910 199150 84980
rect 199350 84910 199360 84980
rect 199140 84860 199360 84910
rect 199640 85090 199860 85140
rect 199640 85020 199650 85090
rect 199850 85020 199860 85090
rect 199640 84980 199860 85020
rect 199640 84910 199650 84980
rect 199850 84910 199860 84980
rect 199640 84860 199860 84910
rect 200140 85090 200360 85140
rect 200140 85020 200150 85090
rect 200350 85020 200360 85090
rect 200140 84980 200360 85020
rect 200140 84910 200150 84980
rect 200350 84910 200360 84980
rect 200140 84860 200360 84910
rect 200640 85090 200860 85140
rect 200640 85020 200650 85090
rect 200850 85020 200860 85090
rect 200640 84980 200860 85020
rect 200640 84910 200650 84980
rect 200850 84910 200860 84980
rect 200640 84860 200860 84910
rect 201140 85090 201360 85140
rect 201140 85020 201150 85090
rect 201350 85020 201360 85090
rect 201140 84980 201360 85020
rect 201140 84910 201150 84980
rect 201350 84910 201360 84980
rect 201140 84860 201360 84910
rect 201640 85090 201860 85140
rect 201640 85020 201650 85090
rect 201850 85020 201860 85090
rect 201640 84980 201860 85020
rect 201640 84910 201650 84980
rect 201850 84910 201860 84980
rect 201640 84860 201860 84910
rect 202140 85090 202360 85140
rect 202140 85020 202150 85090
rect 202350 85020 202360 85090
rect 202140 84980 202360 85020
rect 202140 84910 202150 84980
rect 202350 84910 202360 84980
rect 202140 84860 202360 84910
rect 202640 85090 202860 85140
rect 202640 85020 202650 85090
rect 202850 85020 202860 85090
rect 202640 84980 202860 85020
rect 202640 84910 202650 84980
rect 202850 84910 202860 84980
rect 202640 84860 202860 84910
rect 203140 85090 203360 85140
rect 203140 85020 203150 85090
rect 203350 85020 203360 85090
rect 203140 84980 203360 85020
rect 203140 84910 203150 84980
rect 203350 84910 203360 84980
rect 203140 84860 203360 84910
rect 203640 85090 203860 85140
rect 203640 85020 203650 85090
rect 203850 85020 203860 85090
rect 203640 84980 203860 85020
rect 203640 84910 203650 84980
rect 203850 84910 203860 84980
rect 203640 84860 203860 84910
rect 204140 85090 204360 85140
rect 204140 85020 204150 85090
rect 204350 85020 204360 85090
rect 204140 84980 204360 85020
rect 204140 84910 204150 84980
rect 204350 84910 204360 84980
rect 204140 84860 204360 84910
rect 204640 85090 204860 85140
rect 204640 85020 204650 85090
rect 204850 85020 204860 85090
rect 204640 84980 204860 85020
rect 204640 84910 204650 84980
rect 204850 84910 204860 84980
rect 204640 84860 204860 84910
rect 205140 85090 205360 85140
rect 205140 85020 205150 85090
rect 205350 85020 205360 85090
rect 205140 84980 205360 85020
rect 205140 84910 205150 84980
rect 205350 84910 205360 84980
rect 205140 84860 205360 84910
rect 205640 85090 205860 85140
rect 205640 85020 205650 85090
rect 205850 85020 205860 85090
rect 205640 84980 205860 85020
rect 205640 84910 205650 84980
rect 205850 84910 205860 84980
rect 205640 84860 205860 84910
rect 206140 85090 206360 85140
rect 206140 85020 206150 85090
rect 206350 85020 206360 85090
rect 206140 84980 206360 85020
rect 206140 84910 206150 84980
rect 206350 84910 206360 84980
rect 206140 84860 206360 84910
rect 206640 85090 206860 85140
rect 206640 85020 206650 85090
rect 206850 85020 206860 85090
rect 206640 84980 206860 85020
rect 206640 84910 206650 84980
rect 206850 84910 206860 84980
rect 206640 84860 206860 84910
rect 207140 85090 207360 85140
rect 207140 85020 207150 85090
rect 207350 85020 207360 85090
rect 207140 84980 207360 85020
rect 207140 84910 207150 84980
rect 207350 84910 207360 84980
rect 207140 84860 207360 84910
rect 207640 85090 207860 85140
rect 207640 85020 207650 85090
rect 207850 85020 207860 85090
rect 207640 84980 207860 85020
rect 207640 84910 207650 84980
rect 207850 84910 207860 84980
rect 207640 84860 207860 84910
rect 196000 84850 208000 84860
rect 196000 84650 196020 84850
rect 196090 84650 196410 84850
rect 196480 84650 196520 84850
rect 196590 84650 196910 84850
rect 196980 84650 197020 84850
rect 197090 84650 197410 84850
rect 197480 84650 197520 84850
rect 197590 84650 197910 84850
rect 197980 84650 198020 84850
rect 198090 84650 198410 84850
rect 198480 84650 198520 84850
rect 198590 84650 198910 84850
rect 198980 84650 199020 84850
rect 199090 84650 199410 84850
rect 199480 84650 199520 84850
rect 199590 84650 199910 84850
rect 199980 84650 200020 84850
rect 200090 84650 200410 84850
rect 200480 84650 200520 84850
rect 200590 84650 200910 84850
rect 200980 84650 201020 84850
rect 201090 84650 201410 84850
rect 201480 84650 201520 84850
rect 201590 84650 201910 84850
rect 201980 84650 202020 84850
rect 202090 84650 202410 84850
rect 202480 84650 202520 84850
rect 202590 84650 202910 84850
rect 202980 84650 203020 84850
rect 203090 84650 203410 84850
rect 203480 84650 203520 84850
rect 203590 84650 203910 84850
rect 203980 84650 204020 84850
rect 204090 84650 204410 84850
rect 204480 84650 204520 84850
rect 204590 84650 204910 84850
rect 204980 84650 205020 84850
rect 205090 84650 205410 84850
rect 205480 84650 205520 84850
rect 205590 84650 205910 84850
rect 205980 84650 206020 84850
rect 206090 84650 206410 84850
rect 206480 84650 206520 84850
rect 206590 84650 206910 84850
rect 206980 84650 207020 84850
rect 207090 84650 207410 84850
rect 207480 84650 207520 84850
rect 207590 84650 207910 84850
rect 207980 84650 208000 84850
rect 196000 84640 208000 84650
rect 196140 84590 196360 84640
rect 196140 84520 196150 84590
rect 196350 84520 196360 84590
rect 196140 84480 196360 84520
rect 196140 84410 196150 84480
rect 196350 84410 196360 84480
rect 196140 84360 196360 84410
rect 196640 84590 196860 84640
rect 196640 84520 196650 84590
rect 196850 84520 196860 84590
rect 196640 84480 196860 84520
rect 196640 84410 196650 84480
rect 196850 84410 196860 84480
rect 196640 84360 196860 84410
rect 197140 84590 197360 84640
rect 197140 84520 197150 84590
rect 197350 84520 197360 84590
rect 197140 84480 197360 84520
rect 197140 84410 197150 84480
rect 197350 84410 197360 84480
rect 197140 84360 197360 84410
rect 197640 84590 197860 84640
rect 197640 84520 197650 84590
rect 197850 84520 197860 84590
rect 197640 84480 197860 84520
rect 197640 84410 197650 84480
rect 197850 84410 197860 84480
rect 197640 84360 197860 84410
rect 198140 84590 198360 84640
rect 198140 84520 198150 84590
rect 198350 84520 198360 84590
rect 198140 84480 198360 84520
rect 198140 84410 198150 84480
rect 198350 84410 198360 84480
rect 198140 84360 198360 84410
rect 198640 84590 198860 84640
rect 198640 84520 198650 84590
rect 198850 84520 198860 84590
rect 198640 84480 198860 84520
rect 198640 84410 198650 84480
rect 198850 84410 198860 84480
rect 198640 84360 198860 84410
rect 199140 84590 199360 84640
rect 199140 84520 199150 84590
rect 199350 84520 199360 84590
rect 199140 84480 199360 84520
rect 199140 84410 199150 84480
rect 199350 84410 199360 84480
rect 199140 84360 199360 84410
rect 199640 84590 199860 84640
rect 199640 84520 199650 84590
rect 199850 84520 199860 84590
rect 199640 84480 199860 84520
rect 199640 84410 199650 84480
rect 199850 84410 199860 84480
rect 199640 84360 199860 84410
rect 200140 84590 200360 84640
rect 200140 84520 200150 84590
rect 200350 84520 200360 84590
rect 200140 84480 200360 84520
rect 200140 84410 200150 84480
rect 200350 84410 200360 84480
rect 200140 84360 200360 84410
rect 200640 84590 200860 84640
rect 200640 84520 200650 84590
rect 200850 84520 200860 84590
rect 200640 84480 200860 84520
rect 200640 84410 200650 84480
rect 200850 84410 200860 84480
rect 200640 84360 200860 84410
rect 201140 84590 201360 84640
rect 201140 84520 201150 84590
rect 201350 84520 201360 84590
rect 201140 84480 201360 84520
rect 201140 84410 201150 84480
rect 201350 84410 201360 84480
rect 201140 84360 201360 84410
rect 201640 84590 201860 84640
rect 201640 84520 201650 84590
rect 201850 84520 201860 84590
rect 201640 84480 201860 84520
rect 201640 84410 201650 84480
rect 201850 84410 201860 84480
rect 201640 84360 201860 84410
rect 202140 84590 202360 84640
rect 202140 84520 202150 84590
rect 202350 84520 202360 84590
rect 202140 84480 202360 84520
rect 202140 84410 202150 84480
rect 202350 84410 202360 84480
rect 202140 84360 202360 84410
rect 202640 84590 202860 84640
rect 202640 84520 202650 84590
rect 202850 84520 202860 84590
rect 202640 84480 202860 84520
rect 202640 84410 202650 84480
rect 202850 84410 202860 84480
rect 202640 84360 202860 84410
rect 203140 84590 203360 84640
rect 203140 84520 203150 84590
rect 203350 84520 203360 84590
rect 203140 84480 203360 84520
rect 203140 84410 203150 84480
rect 203350 84410 203360 84480
rect 203140 84360 203360 84410
rect 203640 84590 203860 84640
rect 203640 84520 203650 84590
rect 203850 84520 203860 84590
rect 203640 84480 203860 84520
rect 203640 84410 203650 84480
rect 203850 84410 203860 84480
rect 203640 84360 203860 84410
rect 204140 84590 204360 84640
rect 204140 84520 204150 84590
rect 204350 84520 204360 84590
rect 204140 84480 204360 84520
rect 204140 84410 204150 84480
rect 204350 84410 204360 84480
rect 204140 84360 204360 84410
rect 204640 84590 204860 84640
rect 204640 84520 204650 84590
rect 204850 84520 204860 84590
rect 204640 84480 204860 84520
rect 204640 84410 204650 84480
rect 204850 84410 204860 84480
rect 204640 84360 204860 84410
rect 205140 84590 205360 84640
rect 205140 84520 205150 84590
rect 205350 84520 205360 84590
rect 205140 84480 205360 84520
rect 205140 84410 205150 84480
rect 205350 84410 205360 84480
rect 205140 84360 205360 84410
rect 205640 84590 205860 84640
rect 205640 84520 205650 84590
rect 205850 84520 205860 84590
rect 205640 84480 205860 84520
rect 205640 84410 205650 84480
rect 205850 84410 205860 84480
rect 205640 84360 205860 84410
rect 206140 84590 206360 84640
rect 206140 84520 206150 84590
rect 206350 84520 206360 84590
rect 206140 84480 206360 84520
rect 206140 84410 206150 84480
rect 206350 84410 206360 84480
rect 206140 84360 206360 84410
rect 206640 84590 206860 84640
rect 206640 84520 206650 84590
rect 206850 84520 206860 84590
rect 206640 84480 206860 84520
rect 206640 84410 206650 84480
rect 206850 84410 206860 84480
rect 206640 84360 206860 84410
rect 207140 84590 207360 84640
rect 207140 84520 207150 84590
rect 207350 84520 207360 84590
rect 207140 84480 207360 84520
rect 207140 84410 207150 84480
rect 207350 84410 207360 84480
rect 207140 84360 207360 84410
rect 207640 84590 207860 84640
rect 207640 84520 207650 84590
rect 207850 84520 207860 84590
rect 207640 84480 207860 84520
rect 207640 84410 207650 84480
rect 207850 84410 207860 84480
rect 207640 84360 207860 84410
rect 196000 84350 208000 84360
rect 196000 84150 196020 84350
rect 196090 84150 196410 84350
rect 196480 84150 196520 84350
rect 196590 84150 196910 84350
rect 196980 84150 197020 84350
rect 197090 84150 197410 84350
rect 197480 84150 197520 84350
rect 197590 84150 197910 84350
rect 197980 84150 198020 84350
rect 198090 84150 198410 84350
rect 198480 84150 198520 84350
rect 198590 84150 198910 84350
rect 198980 84150 199020 84350
rect 199090 84150 199410 84350
rect 199480 84150 199520 84350
rect 199590 84150 199910 84350
rect 199980 84150 200020 84350
rect 200090 84150 200410 84350
rect 200480 84150 200520 84350
rect 200590 84150 200910 84350
rect 200980 84150 201020 84350
rect 201090 84150 201410 84350
rect 201480 84150 201520 84350
rect 201590 84150 201910 84350
rect 201980 84150 202020 84350
rect 202090 84150 202410 84350
rect 202480 84150 202520 84350
rect 202590 84150 202910 84350
rect 202980 84150 203020 84350
rect 203090 84150 203410 84350
rect 203480 84150 203520 84350
rect 203590 84150 203910 84350
rect 203980 84150 204020 84350
rect 204090 84150 204410 84350
rect 204480 84150 204520 84350
rect 204590 84150 204910 84350
rect 204980 84150 205020 84350
rect 205090 84150 205410 84350
rect 205480 84150 205520 84350
rect 205590 84150 205910 84350
rect 205980 84150 206020 84350
rect 206090 84150 206410 84350
rect 206480 84150 206520 84350
rect 206590 84150 206910 84350
rect 206980 84150 207020 84350
rect 207090 84150 207410 84350
rect 207480 84150 207520 84350
rect 207590 84150 207910 84350
rect 207980 84150 208000 84350
rect 196000 84140 208000 84150
rect 196140 84090 196360 84140
rect 196140 84020 196150 84090
rect 196350 84020 196360 84090
rect 196140 83980 196360 84020
rect 196140 83910 196150 83980
rect 196350 83910 196360 83980
rect 196140 83860 196360 83910
rect 196640 84090 196860 84140
rect 196640 84020 196650 84090
rect 196850 84020 196860 84090
rect 196640 83980 196860 84020
rect 196640 83910 196650 83980
rect 196850 83910 196860 83980
rect 196640 83860 196860 83910
rect 197140 84090 197360 84140
rect 197140 84020 197150 84090
rect 197350 84020 197360 84090
rect 197140 83980 197360 84020
rect 197140 83910 197150 83980
rect 197350 83910 197360 83980
rect 197140 83860 197360 83910
rect 197640 84090 197860 84140
rect 197640 84020 197650 84090
rect 197850 84020 197860 84090
rect 197640 83980 197860 84020
rect 197640 83910 197650 83980
rect 197850 83910 197860 83980
rect 197640 83860 197860 83910
rect 198140 84090 198360 84140
rect 198140 84020 198150 84090
rect 198350 84020 198360 84090
rect 198140 83980 198360 84020
rect 198140 83910 198150 83980
rect 198350 83910 198360 83980
rect 198140 83860 198360 83910
rect 198640 84090 198860 84140
rect 198640 84020 198650 84090
rect 198850 84020 198860 84090
rect 198640 83980 198860 84020
rect 198640 83910 198650 83980
rect 198850 83910 198860 83980
rect 198640 83860 198860 83910
rect 199140 84090 199360 84140
rect 199140 84020 199150 84090
rect 199350 84020 199360 84090
rect 199140 83980 199360 84020
rect 199140 83910 199150 83980
rect 199350 83910 199360 83980
rect 199140 83860 199360 83910
rect 199640 84090 199860 84140
rect 199640 84020 199650 84090
rect 199850 84020 199860 84090
rect 199640 83980 199860 84020
rect 199640 83910 199650 83980
rect 199850 83910 199860 83980
rect 199640 83860 199860 83910
rect 200140 84090 200360 84140
rect 200140 84020 200150 84090
rect 200350 84020 200360 84090
rect 200140 83980 200360 84020
rect 200140 83910 200150 83980
rect 200350 83910 200360 83980
rect 200140 83860 200360 83910
rect 200640 84090 200860 84140
rect 200640 84020 200650 84090
rect 200850 84020 200860 84090
rect 200640 83980 200860 84020
rect 200640 83910 200650 83980
rect 200850 83910 200860 83980
rect 200640 83860 200860 83910
rect 201140 84090 201360 84140
rect 201140 84020 201150 84090
rect 201350 84020 201360 84090
rect 201140 83980 201360 84020
rect 201140 83910 201150 83980
rect 201350 83910 201360 83980
rect 201140 83860 201360 83910
rect 201640 84090 201860 84140
rect 201640 84020 201650 84090
rect 201850 84020 201860 84090
rect 201640 83980 201860 84020
rect 201640 83910 201650 83980
rect 201850 83910 201860 83980
rect 201640 83860 201860 83910
rect 202140 84090 202360 84140
rect 202140 84020 202150 84090
rect 202350 84020 202360 84090
rect 202140 83980 202360 84020
rect 202140 83910 202150 83980
rect 202350 83910 202360 83980
rect 202140 83860 202360 83910
rect 202640 84090 202860 84140
rect 202640 84020 202650 84090
rect 202850 84020 202860 84090
rect 202640 83980 202860 84020
rect 202640 83910 202650 83980
rect 202850 83910 202860 83980
rect 202640 83860 202860 83910
rect 203140 84090 203360 84140
rect 203140 84020 203150 84090
rect 203350 84020 203360 84090
rect 203140 83980 203360 84020
rect 203140 83910 203150 83980
rect 203350 83910 203360 83980
rect 203140 83860 203360 83910
rect 203640 84090 203860 84140
rect 203640 84020 203650 84090
rect 203850 84020 203860 84090
rect 203640 83980 203860 84020
rect 203640 83910 203650 83980
rect 203850 83910 203860 83980
rect 203640 83860 203860 83910
rect 204140 84090 204360 84140
rect 204140 84020 204150 84090
rect 204350 84020 204360 84090
rect 204140 83980 204360 84020
rect 204140 83910 204150 83980
rect 204350 83910 204360 83980
rect 204140 83860 204360 83910
rect 204640 84090 204860 84140
rect 204640 84020 204650 84090
rect 204850 84020 204860 84090
rect 204640 83980 204860 84020
rect 204640 83910 204650 83980
rect 204850 83910 204860 83980
rect 204640 83860 204860 83910
rect 205140 84090 205360 84140
rect 205140 84020 205150 84090
rect 205350 84020 205360 84090
rect 205140 83980 205360 84020
rect 205140 83910 205150 83980
rect 205350 83910 205360 83980
rect 205140 83860 205360 83910
rect 205640 84090 205860 84140
rect 205640 84020 205650 84090
rect 205850 84020 205860 84090
rect 205640 83980 205860 84020
rect 205640 83910 205650 83980
rect 205850 83910 205860 83980
rect 205640 83860 205860 83910
rect 206140 84090 206360 84140
rect 206140 84020 206150 84090
rect 206350 84020 206360 84090
rect 206140 83980 206360 84020
rect 206140 83910 206150 83980
rect 206350 83910 206360 83980
rect 206140 83860 206360 83910
rect 206640 84090 206860 84140
rect 206640 84020 206650 84090
rect 206850 84020 206860 84090
rect 206640 83980 206860 84020
rect 206640 83910 206650 83980
rect 206850 83910 206860 83980
rect 206640 83860 206860 83910
rect 207140 84090 207360 84140
rect 207140 84020 207150 84090
rect 207350 84020 207360 84090
rect 207140 83980 207360 84020
rect 207140 83910 207150 83980
rect 207350 83910 207360 83980
rect 207140 83860 207360 83910
rect 207640 84090 207860 84140
rect 207640 84020 207650 84090
rect 207850 84020 207860 84090
rect 207640 83980 207860 84020
rect 207640 83910 207650 83980
rect 207850 83910 207860 83980
rect 207640 83860 207860 83910
rect 196000 83850 208000 83860
rect 196000 83650 196020 83850
rect 196090 83650 196410 83850
rect 196480 83650 196520 83850
rect 196590 83650 196910 83850
rect 196980 83650 197020 83850
rect 197090 83650 197410 83850
rect 197480 83650 197520 83850
rect 197590 83650 197910 83850
rect 197980 83650 198020 83850
rect 198090 83650 198410 83850
rect 198480 83650 198520 83850
rect 198590 83650 198910 83850
rect 198980 83650 199020 83850
rect 199090 83650 199410 83850
rect 199480 83650 199520 83850
rect 199590 83650 199910 83850
rect 199980 83650 200020 83850
rect 200090 83650 200410 83850
rect 200480 83650 200520 83850
rect 200590 83650 200910 83850
rect 200980 83650 201020 83850
rect 201090 83650 201410 83850
rect 201480 83650 201520 83850
rect 201590 83650 201910 83850
rect 201980 83650 202020 83850
rect 202090 83650 202410 83850
rect 202480 83650 202520 83850
rect 202590 83650 202910 83850
rect 202980 83650 203020 83850
rect 203090 83650 203410 83850
rect 203480 83650 203520 83850
rect 203590 83650 203910 83850
rect 203980 83650 204020 83850
rect 204090 83650 204410 83850
rect 204480 83650 204520 83850
rect 204590 83650 204910 83850
rect 204980 83650 205020 83850
rect 205090 83650 205410 83850
rect 205480 83650 205520 83850
rect 205590 83650 205910 83850
rect 205980 83650 206020 83850
rect 206090 83650 206410 83850
rect 206480 83650 206520 83850
rect 206590 83650 206910 83850
rect 206980 83650 207020 83850
rect 207090 83650 207410 83850
rect 207480 83650 207520 83850
rect 207590 83650 207910 83850
rect 207980 83650 208000 83850
rect 196000 83640 208000 83650
rect 196140 83590 196360 83640
rect 196140 83520 196150 83590
rect 196350 83520 196360 83590
rect 196140 83480 196360 83520
rect 196140 83410 196150 83480
rect 196350 83410 196360 83480
rect 196140 83360 196360 83410
rect 196640 83590 196860 83640
rect 196640 83520 196650 83590
rect 196850 83520 196860 83590
rect 196640 83480 196860 83520
rect 196640 83410 196650 83480
rect 196850 83410 196860 83480
rect 196640 83360 196860 83410
rect 197140 83590 197360 83640
rect 197140 83520 197150 83590
rect 197350 83520 197360 83590
rect 197140 83480 197360 83520
rect 197140 83410 197150 83480
rect 197350 83410 197360 83480
rect 197140 83360 197360 83410
rect 197640 83590 197860 83640
rect 197640 83520 197650 83590
rect 197850 83520 197860 83590
rect 197640 83480 197860 83520
rect 197640 83410 197650 83480
rect 197850 83410 197860 83480
rect 197640 83360 197860 83410
rect 198140 83590 198360 83640
rect 198140 83520 198150 83590
rect 198350 83520 198360 83590
rect 198140 83480 198360 83520
rect 198140 83410 198150 83480
rect 198350 83410 198360 83480
rect 198140 83360 198360 83410
rect 198640 83590 198860 83640
rect 198640 83520 198650 83590
rect 198850 83520 198860 83590
rect 198640 83480 198860 83520
rect 198640 83410 198650 83480
rect 198850 83410 198860 83480
rect 198640 83360 198860 83410
rect 199140 83590 199360 83640
rect 199140 83520 199150 83590
rect 199350 83520 199360 83590
rect 199140 83480 199360 83520
rect 199140 83410 199150 83480
rect 199350 83410 199360 83480
rect 199140 83360 199360 83410
rect 199640 83590 199860 83640
rect 199640 83520 199650 83590
rect 199850 83520 199860 83590
rect 199640 83480 199860 83520
rect 199640 83410 199650 83480
rect 199850 83410 199860 83480
rect 199640 83360 199860 83410
rect 200140 83590 200360 83640
rect 200140 83520 200150 83590
rect 200350 83520 200360 83590
rect 200140 83480 200360 83520
rect 200140 83410 200150 83480
rect 200350 83410 200360 83480
rect 200140 83360 200360 83410
rect 200640 83590 200860 83640
rect 200640 83520 200650 83590
rect 200850 83520 200860 83590
rect 200640 83480 200860 83520
rect 200640 83410 200650 83480
rect 200850 83410 200860 83480
rect 200640 83360 200860 83410
rect 201140 83590 201360 83640
rect 201140 83520 201150 83590
rect 201350 83520 201360 83590
rect 201140 83480 201360 83520
rect 201140 83410 201150 83480
rect 201350 83410 201360 83480
rect 201140 83360 201360 83410
rect 201640 83590 201860 83640
rect 201640 83520 201650 83590
rect 201850 83520 201860 83590
rect 201640 83480 201860 83520
rect 201640 83410 201650 83480
rect 201850 83410 201860 83480
rect 201640 83360 201860 83410
rect 202140 83590 202360 83640
rect 202140 83520 202150 83590
rect 202350 83520 202360 83590
rect 202140 83480 202360 83520
rect 202140 83410 202150 83480
rect 202350 83410 202360 83480
rect 202140 83360 202360 83410
rect 202640 83590 202860 83640
rect 202640 83520 202650 83590
rect 202850 83520 202860 83590
rect 202640 83480 202860 83520
rect 202640 83410 202650 83480
rect 202850 83410 202860 83480
rect 202640 83360 202860 83410
rect 203140 83590 203360 83640
rect 203140 83520 203150 83590
rect 203350 83520 203360 83590
rect 203140 83480 203360 83520
rect 203140 83410 203150 83480
rect 203350 83410 203360 83480
rect 203140 83360 203360 83410
rect 203640 83590 203860 83640
rect 203640 83520 203650 83590
rect 203850 83520 203860 83590
rect 203640 83480 203860 83520
rect 203640 83410 203650 83480
rect 203850 83410 203860 83480
rect 203640 83360 203860 83410
rect 204140 83590 204360 83640
rect 204140 83520 204150 83590
rect 204350 83520 204360 83590
rect 204140 83480 204360 83520
rect 204140 83410 204150 83480
rect 204350 83410 204360 83480
rect 204140 83360 204360 83410
rect 204640 83590 204860 83640
rect 204640 83520 204650 83590
rect 204850 83520 204860 83590
rect 204640 83480 204860 83520
rect 204640 83410 204650 83480
rect 204850 83410 204860 83480
rect 204640 83360 204860 83410
rect 205140 83590 205360 83640
rect 205140 83520 205150 83590
rect 205350 83520 205360 83590
rect 205140 83480 205360 83520
rect 205140 83410 205150 83480
rect 205350 83410 205360 83480
rect 205140 83360 205360 83410
rect 205640 83590 205860 83640
rect 205640 83520 205650 83590
rect 205850 83520 205860 83590
rect 205640 83480 205860 83520
rect 205640 83410 205650 83480
rect 205850 83410 205860 83480
rect 205640 83360 205860 83410
rect 206140 83590 206360 83640
rect 206140 83520 206150 83590
rect 206350 83520 206360 83590
rect 206140 83480 206360 83520
rect 206140 83410 206150 83480
rect 206350 83410 206360 83480
rect 206140 83360 206360 83410
rect 206640 83590 206860 83640
rect 206640 83520 206650 83590
rect 206850 83520 206860 83590
rect 206640 83480 206860 83520
rect 206640 83410 206650 83480
rect 206850 83410 206860 83480
rect 206640 83360 206860 83410
rect 207140 83590 207360 83640
rect 207140 83520 207150 83590
rect 207350 83520 207360 83590
rect 207140 83480 207360 83520
rect 207140 83410 207150 83480
rect 207350 83410 207360 83480
rect 207140 83360 207360 83410
rect 207640 83590 207860 83640
rect 207640 83520 207650 83590
rect 207850 83520 207860 83590
rect 207640 83480 207860 83520
rect 207640 83410 207650 83480
rect 207850 83410 207860 83480
rect 207640 83360 207860 83410
rect 196000 83350 208000 83360
rect 196000 83150 196020 83350
rect 196090 83150 196410 83350
rect 196480 83150 196520 83350
rect 196590 83150 196910 83350
rect 196980 83150 197020 83350
rect 197090 83150 197410 83350
rect 197480 83150 197520 83350
rect 197590 83150 197910 83350
rect 197980 83150 198020 83350
rect 198090 83150 198410 83350
rect 198480 83150 198520 83350
rect 198590 83150 198910 83350
rect 198980 83150 199020 83350
rect 199090 83150 199410 83350
rect 199480 83150 199520 83350
rect 199590 83150 199910 83350
rect 199980 83150 200020 83350
rect 200090 83150 200410 83350
rect 200480 83150 200520 83350
rect 200590 83150 200910 83350
rect 200980 83150 201020 83350
rect 201090 83150 201410 83350
rect 201480 83150 201520 83350
rect 201590 83150 201910 83350
rect 201980 83150 202020 83350
rect 202090 83150 202410 83350
rect 202480 83150 202520 83350
rect 202590 83150 202910 83350
rect 202980 83150 203020 83350
rect 203090 83150 203410 83350
rect 203480 83150 203520 83350
rect 203590 83150 203910 83350
rect 203980 83150 204020 83350
rect 204090 83150 204410 83350
rect 204480 83150 204520 83350
rect 204590 83150 204910 83350
rect 204980 83150 205020 83350
rect 205090 83150 205410 83350
rect 205480 83150 205520 83350
rect 205590 83150 205910 83350
rect 205980 83150 206020 83350
rect 206090 83150 206410 83350
rect 206480 83150 206520 83350
rect 206590 83150 206910 83350
rect 206980 83150 207020 83350
rect 207090 83150 207410 83350
rect 207480 83150 207520 83350
rect 207590 83150 207910 83350
rect 207980 83150 208000 83350
rect 196000 83140 208000 83150
rect 196140 83090 196360 83140
rect 196140 83020 196150 83090
rect 196350 83020 196360 83090
rect 196140 82980 196360 83020
rect 196140 82910 196150 82980
rect 196350 82910 196360 82980
rect 196140 82860 196360 82910
rect 196640 83090 196860 83140
rect 196640 83020 196650 83090
rect 196850 83020 196860 83090
rect 196640 82980 196860 83020
rect 196640 82910 196650 82980
rect 196850 82910 196860 82980
rect 196640 82860 196860 82910
rect 197140 83090 197360 83140
rect 197140 83020 197150 83090
rect 197350 83020 197360 83090
rect 197140 82980 197360 83020
rect 197140 82910 197150 82980
rect 197350 82910 197360 82980
rect 197140 82860 197360 82910
rect 197640 83090 197860 83140
rect 197640 83020 197650 83090
rect 197850 83020 197860 83090
rect 197640 82980 197860 83020
rect 197640 82910 197650 82980
rect 197850 82910 197860 82980
rect 197640 82860 197860 82910
rect 198140 83090 198360 83140
rect 198140 83020 198150 83090
rect 198350 83020 198360 83090
rect 198140 82980 198360 83020
rect 198140 82910 198150 82980
rect 198350 82910 198360 82980
rect 198140 82860 198360 82910
rect 198640 83090 198860 83140
rect 198640 83020 198650 83090
rect 198850 83020 198860 83090
rect 198640 82980 198860 83020
rect 198640 82910 198650 82980
rect 198850 82910 198860 82980
rect 198640 82860 198860 82910
rect 199140 83090 199360 83140
rect 199140 83020 199150 83090
rect 199350 83020 199360 83090
rect 199140 82980 199360 83020
rect 199140 82910 199150 82980
rect 199350 82910 199360 82980
rect 199140 82860 199360 82910
rect 199640 83090 199860 83140
rect 199640 83020 199650 83090
rect 199850 83020 199860 83090
rect 199640 82980 199860 83020
rect 199640 82910 199650 82980
rect 199850 82910 199860 82980
rect 199640 82860 199860 82910
rect 200140 83090 200360 83140
rect 200140 83020 200150 83090
rect 200350 83020 200360 83090
rect 200140 82980 200360 83020
rect 200140 82910 200150 82980
rect 200350 82910 200360 82980
rect 200140 82860 200360 82910
rect 200640 83090 200860 83140
rect 200640 83020 200650 83090
rect 200850 83020 200860 83090
rect 200640 82980 200860 83020
rect 200640 82910 200650 82980
rect 200850 82910 200860 82980
rect 200640 82860 200860 82910
rect 201140 83090 201360 83140
rect 201140 83020 201150 83090
rect 201350 83020 201360 83090
rect 201140 82980 201360 83020
rect 201140 82910 201150 82980
rect 201350 82910 201360 82980
rect 201140 82860 201360 82910
rect 201640 83090 201860 83140
rect 201640 83020 201650 83090
rect 201850 83020 201860 83090
rect 201640 82980 201860 83020
rect 201640 82910 201650 82980
rect 201850 82910 201860 82980
rect 201640 82860 201860 82910
rect 202140 83090 202360 83140
rect 202140 83020 202150 83090
rect 202350 83020 202360 83090
rect 202140 82980 202360 83020
rect 202140 82910 202150 82980
rect 202350 82910 202360 82980
rect 202140 82860 202360 82910
rect 202640 83090 202860 83140
rect 202640 83020 202650 83090
rect 202850 83020 202860 83090
rect 202640 82980 202860 83020
rect 202640 82910 202650 82980
rect 202850 82910 202860 82980
rect 202640 82860 202860 82910
rect 203140 83090 203360 83140
rect 203140 83020 203150 83090
rect 203350 83020 203360 83090
rect 203140 82980 203360 83020
rect 203140 82910 203150 82980
rect 203350 82910 203360 82980
rect 203140 82860 203360 82910
rect 203640 83090 203860 83140
rect 203640 83020 203650 83090
rect 203850 83020 203860 83090
rect 203640 82980 203860 83020
rect 203640 82910 203650 82980
rect 203850 82910 203860 82980
rect 203640 82860 203860 82910
rect 204140 83090 204360 83140
rect 204140 83020 204150 83090
rect 204350 83020 204360 83090
rect 204140 82980 204360 83020
rect 204140 82910 204150 82980
rect 204350 82910 204360 82980
rect 204140 82860 204360 82910
rect 204640 83090 204860 83140
rect 204640 83020 204650 83090
rect 204850 83020 204860 83090
rect 204640 82980 204860 83020
rect 204640 82910 204650 82980
rect 204850 82910 204860 82980
rect 204640 82860 204860 82910
rect 205140 83090 205360 83140
rect 205140 83020 205150 83090
rect 205350 83020 205360 83090
rect 205140 82980 205360 83020
rect 205140 82910 205150 82980
rect 205350 82910 205360 82980
rect 205140 82860 205360 82910
rect 205640 83090 205860 83140
rect 205640 83020 205650 83090
rect 205850 83020 205860 83090
rect 205640 82980 205860 83020
rect 205640 82910 205650 82980
rect 205850 82910 205860 82980
rect 205640 82860 205860 82910
rect 206140 83090 206360 83140
rect 206140 83020 206150 83090
rect 206350 83020 206360 83090
rect 206140 82980 206360 83020
rect 206140 82910 206150 82980
rect 206350 82910 206360 82980
rect 206140 82860 206360 82910
rect 206640 83090 206860 83140
rect 206640 83020 206650 83090
rect 206850 83020 206860 83090
rect 206640 82980 206860 83020
rect 206640 82910 206650 82980
rect 206850 82910 206860 82980
rect 206640 82860 206860 82910
rect 207140 83090 207360 83140
rect 207140 83020 207150 83090
rect 207350 83020 207360 83090
rect 207140 82980 207360 83020
rect 207140 82910 207150 82980
rect 207350 82910 207360 82980
rect 207140 82860 207360 82910
rect 207640 83090 207860 83140
rect 207640 83020 207650 83090
rect 207850 83020 207860 83090
rect 207640 82980 207860 83020
rect 207640 82910 207650 82980
rect 207850 82910 207860 82980
rect 207640 82860 207860 82910
rect 196000 82850 208000 82860
rect 196000 82650 196020 82850
rect 196090 82650 196410 82850
rect 196480 82650 196520 82850
rect 196590 82650 196910 82850
rect 196980 82650 197020 82850
rect 197090 82650 197410 82850
rect 197480 82650 197520 82850
rect 197590 82650 197910 82850
rect 197980 82650 198020 82850
rect 198090 82650 198410 82850
rect 198480 82650 198520 82850
rect 198590 82650 198910 82850
rect 198980 82650 199020 82850
rect 199090 82650 199410 82850
rect 199480 82650 199520 82850
rect 199590 82650 199910 82850
rect 199980 82650 200020 82850
rect 200090 82650 200410 82850
rect 200480 82650 200520 82850
rect 200590 82650 200910 82850
rect 200980 82650 201020 82850
rect 201090 82650 201410 82850
rect 201480 82650 201520 82850
rect 201590 82650 201910 82850
rect 201980 82650 202020 82850
rect 202090 82650 202410 82850
rect 202480 82650 202520 82850
rect 202590 82650 202910 82850
rect 202980 82650 203020 82850
rect 203090 82650 203410 82850
rect 203480 82650 203520 82850
rect 203590 82650 203910 82850
rect 203980 82650 204020 82850
rect 204090 82650 204410 82850
rect 204480 82650 204520 82850
rect 204590 82650 204910 82850
rect 204980 82650 205020 82850
rect 205090 82650 205410 82850
rect 205480 82650 205520 82850
rect 205590 82650 205910 82850
rect 205980 82650 206020 82850
rect 206090 82650 206410 82850
rect 206480 82650 206520 82850
rect 206590 82650 206910 82850
rect 206980 82650 207020 82850
rect 207090 82650 207410 82850
rect 207480 82650 207520 82850
rect 207590 82650 207910 82850
rect 207980 82650 208000 82850
rect 196000 82640 208000 82650
rect 196140 82590 196360 82640
rect 196140 82520 196150 82590
rect 196350 82520 196360 82590
rect 196140 82480 196360 82520
rect 196140 82410 196150 82480
rect 196350 82410 196360 82480
rect 196140 82360 196360 82410
rect 196640 82590 196860 82640
rect 196640 82520 196650 82590
rect 196850 82520 196860 82590
rect 196640 82480 196860 82520
rect 196640 82410 196650 82480
rect 196850 82410 196860 82480
rect 196640 82360 196860 82410
rect 197140 82590 197360 82640
rect 197140 82520 197150 82590
rect 197350 82520 197360 82590
rect 197140 82480 197360 82520
rect 197140 82410 197150 82480
rect 197350 82410 197360 82480
rect 197140 82360 197360 82410
rect 197640 82590 197860 82640
rect 197640 82520 197650 82590
rect 197850 82520 197860 82590
rect 197640 82480 197860 82520
rect 197640 82410 197650 82480
rect 197850 82410 197860 82480
rect 197640 82360 197860 82410
rect 198140 82590 198360 82640
rect 198140 82520 198150 82590
rect 198350 82520 198360 82590
rect 198140 82480 198360 82520
rect 198140 82410 198150 82480
rect 198350 82410 198360 82480
rect 198140 82360 198360 82410
rect 198640 82590 198860 82640
rect 198640 82520 198650 82590
rect 198850 82520 198860 82590
rect 198640 82480 198860 82520
rect 198640 82410 198650 82480
rect 198850 82410 198860 82480
rect 198640 82360 198860 82410
rect 199140 82590 199360 82640
rect 199140 82520 199150 82590
rect 199350 82520 199360 82590
rect 199140 82480 199360 82520
rect 199140 82410 199150 82480
rect 199350 82410 199360 82480
rect 199140 82360 199360 82410
rect 199640 82590 199860 82640
rect 199640 82520 199650 82590
rect 199850 82520 199860 82590
rect 199640 82480 199860 82520
rect 199640 82410 199650 82480
rect 199850 82410 199860 82480
rect 199640 82360 199860 82410
rect 200140 82590 200360 82640
rect 200140 82520 200150 82590
rect 200350 82520 200360 82590
rect 200140 82480 200360 82520
rect 200140 82410 200150 82480
rect 200350 82410 200360 82480
rect 200140 82360 200360 82410
rect 200640 82590 200860 82640
rect 200640 82520 200650 82590
rect 200850 82520 200860 82590
rect 200640 82480 200860 82520
rect 200640 82410 200650 82480
rect 200850 82410 200860 82480
rect 200640 82360 200860 82410
rect 201140 82590 201360 82640
rect 201140 82520 201150 82590
rect 201350 82520 201360 82590
rect 201140 82480 201360 82520
rect 201140 82410 201150 82480
rect 201350 82410 201360 82480
rect 201140 82360 201360 82410
rect 201640 82590 201860 82640
rect 201640 82520 201650 82590
rect 201850 82520 201860 82590
rect 201640 82480 201860 82520
rect 201640 82410 201650 82480
rect 201850 82410 201860 82480
rect 201640 82360 201860 82410
rect 202140 82590 202360 82640
rect 202140 82520 202150 82590
rect 202350 82520 202360 82590
rect 202140 82480 202360 82520
rect 202140 82410 202150 82480
rect 202350 82410 202360 82480
rect 202140 82360 202360 82410
rect 202640 82590 202860 82640
rect 202640 82520 202650 82590
rect 202850 82520 202860 82590
rect 202640 82480 202860 82520
rect 202640 82410 202650 82480
rect 202850 82410 202860 82480
rect 202640 82360 202860 82410
rect 203140 82590 203360 82640
rect 203140 82520 203150 82590
rect 203350 82520 203360 82590
rect 203140 82480 203360 82520
rect 203140 82410 203150 82480
rect 203350 82410 203360 82480
rect 203140 82360 203360 82410
rect 203640 82590 203860 82640
rect 203640 82520 203650 82590
rect 203850 82520 203860 82590
rect 203640 82480 203860 82520
rect 203640 82410 203650 82480
rect 203850 82410 203860 82480
rect 203640 82360 203860 82410
rect 204140 82590 204360 82640
rect 204140 82520 204150 82590
rect 204350 82520 204360 82590
rect 204140 82480 204360 82520
rect 204140 82410 204150 82480
rect 204350 82410 204360 82480
rect 204140 82360 204360 82410
rect 204640 82590 204860 82640
rect 204640 82520 204650 82590
rect 204850 82520 204860 82590
rect 204640 82480 204860 82520
rect 204640 82410 204650 82480
rect 204850 82410 204860 82480
rect 204640 82360 204860 82410
rect 205140 82590 205360 82640
rect 205140 82520 205150 82590
rect 205350 82520 205360 82590
rect 205140 82480 205360 82520
rect 205140 82410 205150 82480
rect 205350 82410 205360 82480
rect 205140 82360 205360 82410
rect 205640 82590 205860 82640
rect 205640 82520 205650 82590
rect 205850 82520 205860 82590
rect 205640 82480 205860 82520
rect 205640 82410 205650 82480
rect 205850 82410 205860 82480
rect 205640 82360 205860 82410
rect 206140 82590 206360 82640
rect 206140 82520 206150 82590
rect 206350 82520 206360 82590
rect 206140 82480 206360 82520
rect 206140 82410 206150 82480
rect 206350 82410 206360 82480
rect 206140 82360 206360 82410
rect 206640 82590 206860 82640
rect 206640 82520 206650 82590
rect 206850 82520 206860 82590
rect 206640 82480 206860 82520
rect 206640 82410 206650 82480
rect 206850 82410 206860 82480
rect 206640 82360 206860 82410
rect 207140 82590 207360 82640
rect 207140 82520 207150 82590
rect 207350 82520 207360 82590
rect 207140 82480 207360 82520
rect 207140 82410 207150 82480
rect 207350 82410 207360 82480
rect 207140 82360 207360 82410
rect 207640 82590 207860 82640
rect 207640 82520 207650 82590
rect 207850 82520 207860 82590
rect 207640 82480 207860 82520
rect 207640 82410 207650 82480
rect 207850 82410 207860 82480
rect 207640 82360 207860 82410
rect 196000 82350 208000 82360
rect 196000 82150 196020 82350
rect 196090 82150 196410 82350
rect 196480 82150 196520 82350
rect 196590 82150 196910 82350
rect 196980 82150 197020 82350
rect 197090 82150 197410 82350
rect 197480 82150 197520 82350
rect 197590 82150 197910 82350
rect 197980 82150 198020 82350
rect 198090 82150 198410 82350
rect 198480 82150 198520 82350
rect 198590 82150 198910 82350
rect 198980 82150 199020 82350
rect 199090 82150 199410 82350
rect 199480 82150 199520 82350
rect 199590 82150 199910 82350
rect 199980 82150 200020 82350
rect 200090 82150 200410 82350
rect 200480 82150 200520 82350
rect 200590 82150 200910 82350
rect 200980 82150 201020 82350
rect 201090 82150 201410 82350
rect 201480 82150 201520 82350
rect 201590 82150 201910 82350
rect 201980 82150 202020 82350
rect 202090 82150 202410 82350
rect 202480 82150 202520 82350
rect 202590 82150 202910 82350
rect 202980 82150 203020 82350
rect 203090 82150 203410 82350
rect 203480 82150 203520 82350
rect 203590 82150 203910 82350
rect 203980 82150 204020 82350
rect 204090 82150 204410 82350
rect 204480 82150 204520 82350
rect 204590 82150 204910 82350
rect 204980 82150 205020 82350
rect 205090 82150 205410 82350
rect 205480 82150 205520 82350
rect 205590 82150 205910 82350
rect 205980 82150 206020 82350
rect 206090 82150 206410 82350
rect 206480 82150 206520 82350
rect 206590 82150 206910 82350
rect 206980 82150 207020 82350
rect 207090 82150 207410 82350
rect 207480 82150 207520 82350
rect 207590 82150 207910 82350
rect 207980 82150 208000 82350
rect 196000 82140 208000 82150
rect 196140 82090 196360 82140
rect 196140 82020 196150 82090
rect 196350 82020 196360 82090
rect 196140 81980 196360 82020
rect 196140 81910 196150 81980
rect 196350 81910 196360 81980
rect 196140 81860 196360 81910
rect 196640 82090 196860 82140
rect 196640 82020 196650 82090
rect 196850 82020 196860 82090
rect 196640 81980 196860 82020
rect 196640 81910 196650 81980
rect 196850 81910 196860 81980
rect 196640 81860 196860 81910
rect 197140 82090 197360 82140
rect 197140 82020 197150 82090
rect 197350 82020 197360 82090
rect 197140 81980 197360 82020
rect 197140 81910 197150 81980
rect 197350 81910 197360 81980
rect 197140 81860 197360 81910
rect 197640 82090 197860 82140
rect 197640 82020 197650 82090
rect 197850 82020 197860 82090
rect 197640 81980 197860 82020
rect 197640 81910 197650 81980
rect 197850 81910 197860 81980
rect 197640 81860 197860 81910
rect 198140 82090 198360 82140
rect 198140 82020 198150 82090
rect 198350 82020 198360 82090
rect 198140 81980 198360 82020
rect 198140 81910 198150 81980
rect 198350 81910 198360 81980
rect 198140 81860 198360 81910
rect 198640 82090 198860 82140
rect 198640 82020 198650 82090
rect 198850 82020 198860 82090
rect 198640 81980 198860 82020
rect 198640 81910 198650 81980
rect 198850 81910 198860 81980
rect 198640 81860 198860 81910
rect 199140 82090 199360 82140
rect 199140 82020 199150 82090
rect 199350 82020 199360 82090
rect 199140 81980 199360 82020
rect 199140 81910 199150 81980
rect 199350 81910 199360 81980
rect 199140 81860 199360 81910
rect 199640 82090 199860 82140
rect 199640 82020 199650 82090
rect 199850 82020 199860 82090
rect 199640 81980 199860 82020
rect 199640 81910 199650 81980
rect 199850 81910 199860 81980
rect 199640 81860 199860 81910
rect 200140 82090 200360 82140
rect 200140 82020 200150 82090
rect 200350 82020 200360 82090
rect 200140 81980 200360 82020
rect 200140 81910 200150 81980
rect 200350 81910 200360 81980
rect 200140 81860 200360 81910
rect 200640 82090 200860 82140
rect 200640 82020 200650 82090
rect 200850 82020 200860 82090
rect 200640 81980 200860 82020
rect 200640 81910 200650 81980
rect 200850 81910 200860 81980
rect 200640 81860 200860 81910
rect 201140 82090 201360 82140
rect 201140 82020 201150 82090
rect 201350 82020 201360 82090
rect 201140 81980 201360 82020
rect 201140 81910 201150 81980
rect 201350 81910 201360 81980
rect 201140 81860 201360 81910
rect 201640 82090 201860 82140
rect 201640 82020 201650 82090
rect 201850 82020 201860 82090
rect 201640 81980 201860 82020
rect 201640 81910 201650 81980
rect 201850 81910 201860 81980
rect 201640 81860 201860 81910
rect 202140 82090 202360 82140
rect 202140 82020 202150 82090
rect 202350 82020 202360 82090
rect 202140 81980 202360 82020
rect 202140 81910 202150 81980
rect 202350 81910 202360 81980
rect 202140 81860 202360 81910
rect 202640 82090 202860 82140
rect 202640 82020 202650 82090
rect 202850 82020 202860 82090
rect 202640 81980 202860 82020
rect 202640 81910 202650 81980
rect 202850 81910 202860 81980
rect 202640 81860 202860 81910
rect 203140 82090 203360 82140
rect 203140 82020 203150 82090
rect 203350 82020 203360 82090
rect 203140 81980 203360 82020
rect 203140 81910 203150 81980
rect 203350 81910 203360 81980
rect 203140 81860 203360 81910
rect 203640 82090 203860 82140
rect 203640 82020 203650 82090
rect 203850 82020 203860 82090
rect 203640 81980 203860 82020
rect 203640 81910 203650 81980
rect 203850 81910 203860 81980
rect 203640 81860 203860 81910
rect 204140 82090 204360 82140
rect 204140 82020 204150 82090
rect 204350 82020 204360 82090
rect 204140 81980 204360 82020
rect 204140 81910 204150 81980
rect 204350 81910 204360 81980
rect 204140 81860 204360 81910
rect 204640 82090 204860 82140
rect 204640 82020 204650 82090
rect 204850 82020 204860 82090
rect 204640 81980 204860 82020
rect 204640 81910 204650 81980
rect 204850 81910 204860 81980
rect 204640 81860 204860 81910
rect 205140 82090 205360 82140
rect 205140 82020 205150 82090
rect 205350 82020 205360 82090
rect 205140 81980 205360 82020
rect 205140 81910 205150 81980
rect 205350 81910 205360 81980
rect 205140 81860 205360 81910
rect 205640 82090 205860 82140
rect 205640 82020 205650 82090
rect 205850 82020 205860 82090
rect 205640 81980 205860 82020
rect 205640 81910 205650 81980
rect 205850 81910 205860 81980
rect 205640 81860 205860 81910
rect 206140 82090 206360 82140
rect 206140 82020 206150 82090
rect 206350 82020 206360 82090
rect 206140 81980 206360 82020
rect 206140 81910 206150 81980
rect 206350 81910 206360 81980
rect 206140 81860 206360 81910
rect 206640 82090 206860 82140
rect 206640 82020 206650 82090
rect 206850 82020 206860 82090
rect 206640 81980 206860 82020
rect 206640 81910 206650 81980
rect 206850 81910 206860 81980
rect 206640 81860 206860 81910
rect 207140 82090 207360 82140
rect 207140 82020 207150 82090
rect 207350 82020 207360 82090
rect 207140 81980 207360 82020
rect 207140 81910 207150 81980
rect 207350 81910 207360 81980
rect 207140 81860 207360 81910
rect 207640 82090 207860 82140
rect 207640 82020 207650 82090
rect 207850 82020 207860 82090
rect 207640 81980 207860 82020
rect 207640 81910 207650 81980
rect 207850 81910 207860 81980
rect 207640 81860 207860 81910
rect 196000 81850 208000 81860
rect 196000 81650 196020 81850
rect 196090 81650 196410 81850
rect 196480 81650 196520 81850
rect 196590 81650 196910 81850
rect 196980 81650 197020 81850
rect 197090 81650 197410 81850
rect 197480 81650 197520 81850
rect 197590 81650 197910 81850
rect 197980 81650 198020 81850
rect 198090 81650 198410 81850
rect 198480 81650 198520 81850
rect 198590 81650 198910 81850
rect 198980 81650 199020 81850
rect 199090 81650 199410 81850
rect 199480 81650 199520 81850
rect 199590 81650 199910 81850
rect 199980 81650 200020 81850
rect 200090 81650 200410 81850
rect 200480 81650 200520 81850
rect 200590 81650 200910 81850
rect 200980 81650 201020 81850
rect 201090 81650 201410 81850
rect 201480 81650 201520 81850
rect 201590 81650 201910 81850
rect 201980 81650 202020 81850
rect 202090 81650 202410 81850
rect 202480 81650 202520 81850
rect 202590 81650 202910 81850
rect 202980 81650 203020 81850
rect 203090 81650 203410 81850
rect 203480 81650 203520 81850
rect 203590 81650 203910 81850
rect 203980 81650 204020 81850
rect 204090 81650 204410 81850
rect 204480 81650 204520 81850
rect 204590 81650 204910 81850
rect 204980 81650 205020 81850
rect 205090 81650 205410 81850
rect 205480 81650 205520 81850
rect 205590 81650 205910 81850
rect 205980 81650 206020 81850
rect 206090 81650 206410 81850
rect 206480 81650 206520 81850
rect 206590 81650 206910 81850
rect 206980 81650 207020 81850
rect 207090 81650 207410 81850
rect 207480 81650 207520 81850
rect 207590 81650 207910 81850
rect 207980 81650 208000 81850
rect 196000 81640 208000 81650
rect 196140 81590 196360 81640
rect 196140 81520 196150 81590
rect 196350 81520 196360 81590
rect 196140 81480 196360 81520
rect 196140 81410 196150 81480
rect 196350 81410 196360 81480
rect 196140 81360 196360 81410
rect 196640 81590 196860 81640
rect 196640 81520 196650 81590
rect 196850 81520 196860 81590
rect 196640 81480 196860 81520
rect 196640 81410 196650 81480
rect 196850 81410 196860 81480
rect 196640 81360 196860 81410
rect 197140 81590 197360 81640
rect 197140 81520 197150 81590
rect 197350 81520 197360 81590
rect 197140 81480 197360 81520
rect 197140 81410 197150 81480
rect 197350 81410 197360 81480
rect 197140 81360 197360 81410
rect 197640 81590 197860 81640
rect 197640 81520 197650 81590
rect 197850 81520 197860 81590
rect 197640 81480 197860 81520
rect 197640 81410 197650 81480
rect 197850 81410 197860 81480
rect 197640 81360 197860 81410
rect 198140 81590 198360 81640
rect 198140 81520 198150 81590
rect 198350 81520 198360 81590
rect 198140 81480 198360 81520
rect 198140 81410 198150 81480
rect 198350 81410 198360 81480
rect 198140 81360 198360 81410
rect 198640 81590 198860 81640
rect 198640 81520 198650 81590
rect 198850 81520 198860 81590
rect 198640 81480 198860 81520
rect 198640 81410 198650 81480
rect 198850 81410 198860 81480
rect 198640 81360 198860 81410
rect 199140 81590 199360 81640
rect 199140 81520 199150 81590
rect 199350 81520 199360 81590
rect 199140 81480 199360 81520
rect 199140 81410 199150 81480
rect 199350 81410 199360 81480
rect 199140 81360 199360 81410
rect 199640 81590 199860 81640
rect 199640 81520 199650 81590
rect 199850 81520 199860 81590
rect 199640 81480 199860 81520
rect 199640 81410 199650 81480
rect 199850 81410 199860 81480
rect 199640 81360 199860 81410
rect 200140 81590 200360 81640
rect 200140 81520 200150 81590
rect 200350 81520 200360 81590
rect 200140 81480 200360 81520
rect 200140 81410 200150 81480
rect 200350 81410 200360 81480
rect 200140 81360 200360 81410
rect 200640 81590 200860 81640
rect 200640 81520 200650 81590
rect 200850 81520 200860 81590
rect 200640 81480 200860 81520
rect 200640 81410 200650 81480
rect 200850 81410 200860 81480
rect 200640 81360 200860 81410
rect 201140 81590 201360 81640
rect 201140 81520 201150 81590
rect 201350 81520 201360 81590
rect 201140 81480 201360 81520
rect 201140 81410 201150 81480
rect 201350 81410 201360 81480
rect 201140 81360 201360 81410
rect 201640 81590 201860 81640
rect 201640 81520 201650 81590
rect 201850 81520 201860 81590
rect 201640 81480 201860 81520
rect 201640 81410 201650 81480
rect 201850 81410 201860 81480
rect 201640 81360 201860 81410
rect 202140 81590 202360 81640
rect 202140 81520 202150 81590
rect 202350 81520 202360 81590
rect 202140 81480 202360 81520
rect 202140 81410 202150 81480
rect 202350 81410 202360 81480
rect 202140 81360 202360 81410
rect 202640 81590 202860 81640
rect 202640 81520 202650 81590
rect 202850 81520 202860 81590
rect 202640 81480 202860 81520
rect 202640 81410 202650 81480
rect 202850 81410 202860 81480
rect 202640 81360 202860 81410
rect 203140 81590 203360 81640
rect 203140 81520 203150 81590
rect 203350 81520 203360 81590
rect 203140 81480 203360 81520
rect 203140 81410 203150 81480
rect 203350 81410 203360 81480
rect 203140 81360 203360 81410
rect 203640 81590 203860 81640
rect 203640 81520 203650 81590
rect 203850 81520 203860 81590
rect 203640 81480 203860 81520
rect 203640 81410 203650 81480
rect 203850 81410 203860 81480
rect 203640 81360 203860 81410
rect 204140 81590 204360 81640
rect 204140 81520 204150 81590
rect 204350 81520 204360 81590
rect 204140 81480 204360 81520
rect 204140 81410 204150 81480
rect 204350 81410 204360 81480
rect 204140 81360 204360 81410
rect 204640 81590 204860 81640
rect 204640 81520 204650 81590
rect 204850 81520 204860 81590
rect 204640 81480 204860 81520
rect 204640 81410 204650 81480
rect 204850 81410 204860 81480
rect 204640 81360 204860 81410
rect 205140 81590 205360 81640
rect 205140 81520 205150 81590
rect 205350 81520 205360 81590
rect 205140 81480 205360 81520
rect 205140 81410 205150 81480
rect 205350 81410 205360 81480
rect 205140 81360 205360 81410
rect 205640 81590 205860 81640
rect 205640 81520 205650 81590
rect 205850 81520 205860 81590
rect 205640 81480 205860 81520
rect 205640 81410 205650 81480
rect 205850 81410 205860 81480
rect 205640 81360 205860 81410
rect 206140 81590 206360 81640
rect 206140 81520 206150 81590
rect 206350 81520 206360 81590
rect 206140 81480 206360 81520
rect 206140 81410 206150 81480
rect 206350 81410 206360 81480
rect 206140 81360 206360 81410
rect 206640 81590 206860 81640
rect 206640 81520 206650 81590
rect 206850 81520 206860 81590
rect 206640 81480 206860 81520
rect 206640 81410 206650 81480
rect 206850 81410 206860 81480
rect 206640 81360 206860 81410
rect 207140 81590 207360 81640
rect 207140 81520 207150 81590
rect 207350 81520 207360 81590
rect 207140 81480 207360 81520
rect 207140 81410 207150 81480
rect 207350 81410 207360 81480
rect 207140 81360 207360 81410
rect 207640 81590 207860 81640
rect 207640 81520 207650 81590
rect 207850 81520 207860 81590
rect 207640 81480 207860 81520
rect 207640 81410 207650 81480
rect 207850 81410 207860 81480
rect 207640 81360 207860 81410
rect 196000 81350 208000 81360
rect 196000 81150 196020 81350
rect 196090 81150 196410 81350
rect 196480 81150 196520 81350
rect 196590 81150 196910 81350
rect 196980 81150 197020 81350
rect 197090 81150 197410 81350
rect 197480 81150 197520 81350
rect 197590 81150 197910 81350
rect 197980 81150 198020 81350
rect 198090 81150 198410 81350
rect 198480 81150 198520 81350
rect 198590 81150 198910 81350
rect 198980 81150 199020 81350
rect 199090 81150 199410 81350
rect 199480 81150 199520 81350
rect 199590 81150 199910 81350
rect 199980 81150 200020 81350
rect 200090 81150 200410 81350
rect 200480 81150 200520 81350
rect 200590 81150 200910 81350
rect 200980 81150 201020 81350
rect 201090 81150 201410 81350
rect 201480 81150 201520 81350
rect 201590 81150 201910 81350
rect 201980 81150 202020 81350
rect 202090 81150 202410 81350
rect 202480 81150 202520 81350
rect 202590 81150 202910 81350
rect 202980 81150 203020 81350
rect 203090 81150 203410 81350
rect 203480 81150 203520 81350
rect 203590 81150 203910 81350
rect 203980 81150 204020 81350
rect 204090 81150 204410 81350
rect 204480 81150 204520 81350
rect 204590 81150 204910 81350
rect 204980 81150 205020 81350
rect 205090 81150 205410 81350
rect 205480 81150 205520 81350
rect 205590 81150 205910 81350
rect 205980 81150 206020 81350
rect 206090 81150 206410 81350
rect 206480 81150 206520 81350
rect 206590 81150 206910 81350
rect 206980 81150 207020 81350
rect 207090 81150 207410 81350
rect 207480 81150 207520 81350
rect 207590 81150 207910 81350
rect 207980 81150 208000 81350
rect 196000 81140 208000 81150
rect 196140 81090 196360 81140
rect 196140 81020 196150 81090
rect 196350 81020 196360 81090
rect 196140 80980 196360 81020
rect 196140 80910 196150 80980
rect 196350 80910 196360 80980
rect 196140 80860 196360 80910
rect 196640 81090 196860 81140
rect 196640 81020 196650 81090
rect 196850 81020 196860 81090
rect 196640 80980 196860 81020
rect 196640 80910 196650 80980
rect 196850 80910 196860 80980
rect 196640 80860 196860 80910
rect 197140 81090 197360 81140
rect 197140 81020 197150 81090
rect 197350 81020 197360 81090
rect 197140 80980 197360 81020
rect 197140 80910 197150 80980
rect 197350 80910 197360 80980
rect 197140 80860 197360 80910
rect 197640 81090 197860 81140
rect 197640 81020 197650 81090
rect 197850 81020 197860 81090
rect 197640 80980 197860 81020
rect 197640 80910 197650 80980
rect 197850 80910 197860 80980
rect 197640 80860 197860 80910
rect 198140 81090 198360 81140
rect 198140 81020 198150 81090
rect 198350 81020 198360 81090
rect 198140 80980 198360 81020
rect 198140 80910 198150 80980
rect 198350 80910 198360 80980
rect 198140 80860 198360 80910
rect 198640 81090 198860 81140
rect 198640 81020 198650 81090
rect 198850 81020 198860 81090
rect 198640 80980 198860 81020
rect 198640 80910 198650 80980
rect 198850 80910 198860 80980
rect 198640 80860 198860 80910
rect 199140 81090 199360 81140
rect 199140 81020 199150 81090
rect 199350 81020 199360 81090
rect 199140 80980 199360 81020
rect 199140 80910 199150 80980
rect 199350 80910 199360 80980
rect 199140 80860 199360 80910
rect 199640 81090 199860 81140
rect 199640 81020 199650 81090
rect 199850 81020 199860 81090
rect 199640 80980 199860 81020
rect 199640 80910 199650 80980
rect 199850 80910 199860 80980
rect 199640 80860 199860 80910
rect 200140 81090 200360 81140
rect 200140 81020 200150 81090
rect 200350 81020 200360 81090
rect 200140 80980 200360 81020
rect 200140 80910 200150 80980
rect 200350 80910 200360 80980
rect 200140 80860 200360 80910
rect 200640 81090 200860 81140
rect 200640 81020 200650 81090
rect 200850 81020 200860 81090
rect 200640 80980 200860 81020
rect 200640 80910 200650 80980
rect 200850 80910 200860 80980
rect 200640 80860 200860 80910
rect 201140 81090 201360 81140
rect 201140 81020 201150 81090
rect 201350 81020 201360 81090
rect 201140 80980 201360 81020
rect 201140 80910 201150 80980
rect 201350 80910 201360 80980
rect 201140 80860 201360 80910
rect 201640 81090 201860 81140
rect 201640 81020 201650 81090
rect 201850 81020 201860 81090
rect 201640 80980 201860 81020
rect 201640 80910 201650 80980
rect 201850 80910 201860 80980
rect 201640 80860 201860 80910
rect 202140 81090 202360 81140
rect 202140 81020 202150 81090
rect 202350 81020 202360 81090
rect 202140 80980 202360 81020
rect 202140 80910 202150 80980
rect 202350 80910 202360 80980
rect 202140 80860 202360 80910
rect 202640 81090 202860 81140
rect 202640 81020 202650 81090
rect 202850 81020 202860 81090
rect 202640 80980 202860 81020
rect 202640 80910 202650 80980
rect 202850 80910 202860 80980
rect 202640 80860 202860 80910
rect 203140 81090 203360 81140
rect 203140 81020 203150 81090
rect 203350 81020 203360 81090
rect 203140 80980 203360 81020
rect 203140 80910 203150 80980
rect 203350 80910 203360 80980
rect 203140 80860 203360 80910
rect 203640 81090 203860 81140
rect 203640 81020 203650 81090
rect 203850 81020 203860 81090
rect 203640 80980 203860 81020
rect 203640 80910 203650 80980
rect 203850 80910 203860 80980
rect 203640 80860 203860 80910
rect 204140 81090 204360 81140
rect 204140 81020 204150 81090
rect 204350 81020 204360 81090
rect 204140 80980 204360 81020
rect 204140 80910 204150 80980
rect 204350 80910 204360 80980
rect 204140 80860 204360 80910
rect 204640 81090 204860 81140
rect 204640 81020 204650 81090
rect 204850 81020 204860 81090
rect 204640 80980 204860 81020
rect 204640 80910 204650 80980
rect 204850 80910 204860 80980
rect 204640 80860 204860 80910
rect 205140 81090 205360 81140
rect 205140 81020 205150 81090
rect 205350 81020 205360 81090
rect 205140 80980 205360 81020
rect 205140 80910 205150 80980
rect 205350 80910 205360 80980
rect 205140 80860 205360 80910
rect 205640 81090 205860 81140
rect 205640 81020 205650 81090
rect 205850 81020 205860 81090
rect 205640 80980 205860 81020
rect 205640 80910 205650 80980
rect 205850 80910 205860 80980
rect 205640 80860 205860 80910
rect 206140 81090 206360 81140
rect 206140 81020 206150 81090
rect 206350 81020 206360 81090
rect 206140 80980 206360 81020
rect 206140 80910 206150 80980
rect 206350 80910 206360 80980
rect 206140 80860 206360 80910
rect 206640 81090 206860 81140
rect 206640 81020 206650 81090
rect 206850 81020 206860 81090
rect 206640 80980 206860 81020
rect 206640 80910 206650 80980
rect 206850 80910 206860 80980
rect 206640 80860 206860 80910
rect 207140 81090 207360 81140
rect 207140 81020 207150 81090
rect 207350 81020 207360 81090
rect 207140 80980 207360 81020
rect 207140 80910 207150 80980
rect 207350 80910 207360 80980
rect 207140 80860 207360 80910
rect 207640 81090 207860 81140
rect 207640 81020 207650 81090
rect 207850 81020 207860 81090
rect 207640 80980 207860 81020
rect 207640 80910 207650 80980
rect 207850 80910 207860 80980
rect 207640 80860 207860 80910
rect 196000 80850 208000 80860
rect 196000 80650 196020 80850
rect 196090 80650 196410 80850
rect 196480 80650 196520 80850
rect 196590 80650 196910 80850
rect 196980 80650 197020 80850
rect 197090 80650 197410 80850
rect 197480 80650 197520 80850
rect 197590 80650 197910 80850
rect 197980 80650 198020 80850
rect 198090 80650 198410 80850
rect 198480 80650 198520 80850
rect 198590 80650 198910 80850
rect 198980 80650 199020 80850
rect 199090 80650 199410 80850
rect 199480 80650 199520 80850
rect 199590 80650 199910 80850
rect 199980 80650 200020 80850
rect 200090 80650 200410 80850
rect 200480 80650 200520 80850
rect 200590 80650 200910 80850
rect 200980 80650 201020 80850
rect 201090 80650 201410 80850
rect 201480 80650 201520 80850
rect 201590 80650 201910 80850
rect 201980 80650 202020 80850
rect 202090 80650 202410 80850
rect 202480 80650 202520 80850
rect 202590 80650 202910 80850
rect 202980 80650 203020 80850
rect 203090 80650 203410 80850
rect 203480 80650 203520 80850
rect 203590 80650 203910 80850
rect 203980 80650 204020 80850
rect 204090 80650 204410 80850
rect 204480 80650 204520 80850
rect 204590 80650 204910 80850
rect 204980 80650 205020 80850
rect 205090 80650 205410 80850
rect 205480 80650 205520 80850
rect 205590 80650 205910 80850
rect 205980 80650 206020 80850
rect 206090 80650 206410 80850
rect 206480 80650 206520 80850
rect 206590 80650 206910 80850
rect 206980 80650 207020 80850
rect 207090 80650 207410 80850
rect 207480 80650 207520 80850
rect 207590 80650 207910 80850
rect 207980 80650 208000 80850
rect 196000 80640 208000 80650
rect 196140 80590 196360 80640
rect 196140 80520 196150 80590
rect 196350 80520 196360 80590
rect 196140 80480 196360 80520
rect 196140 80410 196150 80480
rect 196350 80410 196360 80480
rect 196140 80360 196360 80410
rect 196640 80590 196860 80640
rect 196640 80520 196650 80590
rect 196850 80520 196860 80590
rect 196640 80480 196860 80520
rect 196640 80410 196650 80480
rect 196850 80410 196860 80480
rect 196640 80360 196860 80410
rect 197140 80590 197360 80640
rect 197140 80520 197150 80590
rect 197350 80520 197360 80590
rect 197140 80480 197360 80520
rect 197140 80410 197150 80480
rect 197350 80410 197360 80480
rect 197140 80360 197360 80410
rect 197640 80590 197860 80640
rect 197640 80520 197650 80590
rect 197850 80520 197860 80590
rect 197640 80480 197860 80520
rect 197640 80410 197650 80480
rect 197850 80410 197860 80480
rect 197640 80360 197860 80410
rect 198140 80590 198360 80640
rect 198140 80520 198150 80590
rect 198350 80520 198360 80590
rect 198140 80480 198360 80520
rect 198140 80410 198150 80480
rect 198350 80410 198360 80480
rect 198140 80360 198360 80410
rect 198640 80590 198860 80640
rect 198640 80520 198650 80590
rect 198850 80520 198860 80590
rect 198640 80480 198860 80520
rect 198640 80410 198650 80480
rect 198850 80410 198860 80480
rect 198640 80360 198860 80410
rect 199140 80590 199360 80640
rect 199140 80520 199150 80590
rect 199350 80520 199360 80590
rect 199140 80480 199360 80520
rect 199140 80410 199150 80480
rect 199350 80410 199360 80480
rect 199140 80360 199360 80410
rect 199640 80590 199860 80640
rect 199640 80520 199650 80590
rect 199850 80520 199860 80590
rect 199640 80480 199860 80520
rect 199640 80410 199650 80480
rect 199850 80410 199860 80480
rect 199640 80360 199860 80410
rect 200140 80590 200360 80640
rect 200140 80520 200150 80590
rect 200350 80520 200360 80590
rect 200140 80480 200360 80520
rect 200140 80410 200150 80480
rect 200350 80410 200360 80480
rect 200140 80360 200360 80410
rect 200640 80590 200860 80640
rect 200640 80520 200650 80590
rect 200850 80520 200860 80590
rect 200640 80480 200860 80520
rect 200640 80410 200650 80480
rect 200850 80410 200860 80480
rect 200640 80360 200860 80410
rect 201140 80590 201360 80640
rect 201140 80520 201150 80590
rect 201350 80520 201360 80590
rect 201140 80480 201360 80520
rect 201140 80410 201150 80480
rect 201350 80410 201360 80480
rect 201140 80360 201360 80410
rect 201640 80590 201860 80640
rect 201640 80520 201650 80590
rect 201850 80520 201860 80590
rect 201640 80480 201860 80520
rect 201640 80410 201650 80480
rect 201850 80410 201860 80480
rect 201640 80360 201860 80410
rect 202140 80590 202360 80640
rect 202140 80520 202150 80590
rect 202350 80520 202360 80590
rect 202140 80480 202360 80520
rect 202140 80410 202150 80480
rect 202350 80410 202360 80480
rect 202140 80360 202360 80410
rect 202640 80590 202860 80640
rect 202640 80520 202650 80590
rect 202850 80520 202860 80590
rect 202640 80480 202860 80520
rect 202640 80410 202650 80480
rect 202850 80410 202860 80480
rect 202640 80360 202860 80410
rect 203140 80590 203360 80640
rect 203140 80520 203150 80590
rect 203350 80520 203360 80590
rect 203140 80480 203360 80520
rect 203140 80410 203150 80480
rect 203350 80410 203360 80480
rect 203140 80360 203360 80410
rect 203640 80590 203860 80640
rect 203640 80520 203650 80590
rect 203850 80520 203860 80590
rect 203640 80480 203860 80520
rect 203640 80410 203650 80480
rect 203850 80410 203860 80480
rect 203640 80360 203860 80410
rect 204140 80590 204360 80640
rect 204140 80520 204150 80590
rect 204350 80520 204360 80590
rect 204140 80480 204360 80520
rect 204140 80410 204150 80480
rect 204350 80410 204360 80480
rect 204140 80360 204360 80410
rect 204640 80590 204860 80640
rect 204640 80520 204650 80590
rect 204850 80520 204860 80590
rect 204640 80480 204860 80520
rect 204640 80410 204650 80480
rect 204850 80410 204860 80480
rect 204640 80360 204860 80410
rect 205140 80590 205360 80640
rect 205140 80520 205150 80590
rect 205350 80520 205360 80590
rect 205140 80480 205360 80520
rect 205140 80410 205150 80480
rect 205350 80410 205360 80480
rect 205140 80360 205360 80410
rect 205640 80590 205860 80640
rect 205640 80520 205650 80590
rect 205850 80520 205860 80590
rect 205640 80480 205860 80520
rect 205640 80410 205650 80480
rect 205850 80410 205860 80480
rect 205640 80360 205860 80410
rect 206140 80590 206360 80640
rect 206140 80520 206150 80590
rect 206350 80520 206360 80590
rect 206140 80480 206360 80520
rect 206140 80410 206150 80480
rect 206350 80410 206360 80480
rect 206140 80360 206360 80410
rect 206640 80590 206860 80640
rect 206640 80520 206650 80590
rect 206850 80520 206860 80590
rect 206640 80480 206860 80520
rect 206640 80410 206650 80480
rect 206850 80410 206860 80480
rect 206640 80360 206860 80410
rect 207140 80590 207360 80640
rect 207140 80520 207150 80590
rect 207350 80520 207360 80590
rect 207140 80480 207360 80520
rect 207140 80410 207150 80480
rect 207350 80410 207360 80480
rect 207140 80360 207360 80410
rect 207640 80590 207860 80640
rect 207640 80520 207650 80590
rect 207850 80520 207860 80590
rect 207640 80480 207860 80520
rect 207640 80410 207650 80480
rect 207850 80410 207860 80480
rect 207640 80360 207860 80410
rect 196000 80350 208000 80360
rect 196000 80150 196020 80350
rect 196090 80150 196410 80350
rect 196480 80150 196520 80350
rect 196590 80150 196910 80350
rect 196980 80150 197020 80350
rect 197090 80150 197410 80350
rect 197480 80150 197520 80350
rect 197590 80150 197910 80350
rect 197980 80150 198020 80350
rect 198090 80150 198410 80350
rect 198480 80150 198520 80350
rect 198590 80150 198910 80350
rect 198980 80150 199020 80350
rect 199090 80150 199410 80350
rect 199480 80150 199520 80350
rect 199590 80150 199910 80350
rect 199980 80150 200020 80350
rect 200090 80150 200410 80350
rect 200480 80150 200520 80350
rect 200590 80150 200910 80350
rect 200980 80150 201020 80350
rect 201090 80150 201410 80350
rect 201480 80150 201520 80350
rect 201590 80150 201910 80350
rect 201980 80150 202020 80350
rect 202090 80150 202410 80350
rect 202480 80150 202520 80350
rect 202590 80150 202910 80350
rect 202980 80150 203020 80350
rect 203090 80150 203410 80350
rect 203480 80150 203520 80350
rect 203590 80150 203910 80350
rect 203980 80150 204020 80350
rect 204090 80150 204410 80350
rect 204480 80150 204520 80350
rect 204590 80150 204910 80350
rect 204980 80150 205020 80350
rect 205090 80150 205410 80350
rect 205480 80150 205520 80350
rect 205590 80150 205910 80350
rect 205980 80150 206020 80350
rect 206090 80150 206410 80350
rect 206480 80150 206520 80350
rect 206590 80150 206910 80350
rect 206980 80150 207020 80350
rect 207090 80150 207410 80350
rect 207480 80150 207520 80350
rect 207590 80150 207910 80350
rect 207980 80150 208000 80350
rect 196000 80140 208000 80150
rect 196140 80090 196360 80140
rect 196140 80020 196150 80090
rect 196350 80020 196360 80090
rect 196140 79980 196360 80020
rect 196140 79910 196150 79980
rect 196350 79910 196360 79980
rect 196140 79860 196360 79910
rect 196640 80090 196860 80140
rect 196640 80020 196650 80090
rect 196850 80020 196860 80090
rect 196640 79980 196860 80020
rect 196640 79910 196650 79980
rect 196850 79910 196860 79980
rect 196640 79860 196860 79910
rect 197140 80090 197360 80140
rect 197140 80020 197150 80090
rect 197350 80020 197360 80090
rect 197140 79980 197360 80020
rect 197140 79910 197150 79980
rect 197350 79910 197360 79980
rect 197140 79860 197360 79910
rect 197640 80090 197860 80140
rect 197640 80020 197650 80090
rect 197850 80020 197860 80090
rect 197640 79980 197860 80020
rect 197640 79910 197650 79980
rect 197850 79910 197860 79980
rect 197640 79860 197860 79910
rect 198140 80090 198360 80140
rect 198140 80020 198150 80090
rect 198350 80020 198360 80090
rect 198140 79980 198360 80020
rect 198140 79910 198150 79980
rect 198350 79910 198360 79980
rect 198140 79860 198360 79910
rect 198640 80090 198860 80140
rect 198640 80020 198650 80090
rect 198850 80020 198860 80090
rect 198640 79980 198860 80020
rect 198640 79910 198650 79980
rect 198850 79910 198860 79980
rect 198640 79860 198860 79910
rect 199140 80090 199360 80140
rect 199140 80020 199150 80090
rect 199350 80020 199360 80090
rect 199140 79980 199360 80020
rect 199140 79910 199150 79980
rect 199350 79910 199360 79980
rect 199140 79860 199360 79910
rect 199640 80090 199860 80140
rect 199640 80020 199650 80090
rect 199850 80020 199860 80090
rect 199640 79980 199860 80020
rect 199640 79910 199650 79980
rect 199850 79910 199860 79980
rect 199640 79860 199860 79910
rect 200140 80090 200360 80140
rect 200140 80020 200150 80090
rect 200350 80020 200360 80090
rect 200140 79980 200360 80020
rect 200140 79910 200150 79980
rect 200350 79910 200360 79980
rect 200140 79860 200360 79910
rect 200640 80090 200860 80140
rect 200640 80020 200650 80090
rect 200850 80020 200860 80090
rect 200640 79980 200860 80020
rect 200640 79910 200650 79980
rect 200850 79910 200860 79980
rect 200640 79860 200860 79910
rect 201140 80090 201360 80140
rect 201140 80020 201150 80090
rect 201350 80020 201360 80090
rect 201140 79980 201360 80020
rect 201140 79910 201150 79980
rect 201350 79910 201360 79980
rect 201140 79860 201360 79910
rect 201640 80090 201860 80140
rect 201640 80020 201650 80090
rect 201850 80020 201860 80090
rect 201640 79980 201860 80020
rect 201640 79910 201650 79980
rect 201850 79910 201860 79980
rect 201640 79860 201860 79910
rect 202140 80090 202360 80140
rect 202140 80020 202150 80090
rect 202350 80020 202360 80090
rect 202140 79980 202360 80020
rect 202140 79910 202150 79980
rect 202350 79910 202360 79980
rect 202140 79860 202360 79910
rect 202640 80090 202860 80140
rect 202640 80020 202650 80090
rect 202850 80020 202860 80090
rect 202640 79980 202860 80020
rect 202640 79910 202650 79980
rect 202850 79910 202860 79980
rect 202640 79860 202860 79910
rect 203140 80090 203360 80140
rect 203140 80020 203150 80090
rect 203350 80020 203360 80090
rect 203140 79980 203360 80020
rect 203140 79910 203150 79980
rect 203350 79910 203360 79980
rect 203140 79860 203360 79910
rect 203640 80090 203860 80140
rect 203640 80020 203650 80090
rect 203850 80020 203860 80090
rect 203640 79980 203860 80020
rect 203640 79910 203650 79980
rect 203850 79910 203860 79980
rect 203640 79860 203860 79910
rect 204140 80090 204360 80140
rect 204140 80020 204150 80090
rect 204350 80020 204360 80090
rect 204140 79980 204360 80020
rect 204140 79910 204150 79980
rect 204350 79910 204360 79980
rect 204140 79860 204360 79910
rect 204640 80090 204860 80140
rect 204640 80020 204650 80090
rect 204850 80020 204860 80090
rect 204640 79980 204860 80020
rect 204640 79910 204650 79980
rect 204850 79910 204860 79980
rect 204640 79860 204860 79910
rect 205140 80090 205360 80140
rect 205140 80020 205150 80090
rect 205350 80020 205360 80090
rect 205140 79980 205360 80020
rect 205140 79910 205150 79980
rect 205350 79910 205360 79980
rect 205140 79860 205360 79910
rect 205640 80090 205860 80140
rect 205640 80020 205650 80090
rect 205850 80020 205860 80090
rect 205640 79980 205860 80020
rect 205640 79910 205650 79980
rect 205850 79910 205860 79980
rect 205640 79860 205860 79910
rect 206140 80090 206360 80140
rect 206140 80020 206150 80090
rect 206350 80020 206360 80090
rect 206140 79980 206360 80020
rect 206140 79910 206150 79980
rect 206350 79910 206360 79980
rect 206140 79860 206360 79910
rect 206640 80090 206860 80140
rect 206640 80020 206650 80090
rect 206850 80020 206860 80090
rect 206640 79980 206860 80020
rect 206640 79910 206650 79980
rect 206850 79910 206860 79980
rect 206640 79860 206860 79910
rect 207140 80090 207360 80140
rect 207140 80020 207150 80090
rect 207350 80020 207360 80090
rect 207140 79980 207360 80020
rect 207140 79910 207150 79980
rect 207350 79910 207360 79980
rect 207140 79860 207360 79910
rect 207640 80090 207860 80140
rect 207640 80020 207650 80090
rect 207850 80020 207860 80090
rect 207640 79980 207860 80020
rect 207640 79910 207650 79980
rect 207850 79910 207860 79980
rect 207640 79860 207860 79910
rect 196000 79850 208000 79860
rect 196000 79650 196020 79850
rect 196090 79650 196410 79850
rect 196480 79650 196520 79850
rect 196590 79650 196910 79850
rect 196980 79650 197020 79850
rect 197090 79650 197410 79850
rect 197480 79650 197520 79850
rect 197590 79650 197910 79850
rect 197980 79650 198020 79850
rect 198090 79650 198410 79850
rect 198480 79650 198520 79850
rect 198590 79650 198910 79850
rect 198980 79650 199020 79850
rect 199090 79650 199410 79850
rect 199480 79650 199520 79850
rect 199590 79650 199910 79850
rect 199980 79650 200020 79850
rect 200090 79650 200410 79850
rect 200480 79650 200520 79850
rect 200590 79650 200910 79850
rect 200980 79650 201020 79850
rect 201090 79650 201410 79850
rect 201480 79650 201520 79850
rect 201590 79650 201910 79850
rect 201980 79650 202020 79850
rect 202090 79650 202410 79850
rect 202480 79650 202520 79850
rect 202590 79650 202910 79850
rect 202980 79650 203020 79850
rect 203090 79650 203410 79850
rect 203480 79650 203520 79850
rect 203590 79650 203910 79850
rect 203980 79650 204020 79850
rect 204090 79650 204410 79850
rect 204480 79650 204520 79850
rect 204590 79650 204910 79850
rect 204980 79650 205020 79850
rect 205090 79650 205410 79850
rect 205480 79650 205520 79850
rect 205590 79650 205910 79850
rect 205980 79650 206020 79850
rect 206090 79650 206410 79850
rect 206480 79650 206520 79850
rect 206590 79650 206910 79850
rect 206980 79650 207020 79850
rect 207090 79650 207410 79850
rect 207480 79650 207520 79850
rect 207590 79650 207910 79850
rect 207980 79650 208000 79850
rect 196000 79640 208000 79650
rect 196140 79590 196360 79640
rect 196140 79520 196150 79590
rect 196350 79520 196360 79590
rect 196140 79480 196360 79520
rect 196140 79410 196150 79480
rect 196350 79410 196360 79480
rect 196140 79360 196360 79410
rect 196640 79590 196860 79640
rect 196640 79520 196650 79590
rect 196850 79520 196860 79590
rect 196640 79480 196860 79520
rect 196640 79410 196650 79480
rect 196850 79410 196860 79480
rect 196640 79360 196860 79410
rect 197140 79590 197360 79640
rect 197140 79520 197150 79590
rect 197350 79520 197360 79590
rect 197140 79480 197360 79520
rect 197140 79410 197150 79480
rect 197350 79410 197360 79480
rect 197140 79360 197360 79410
rect 197640 79590 197860 79640
rect 197640 79520 197650 79590
rect 197850 79520 197860 79590
rect 197640 79480 197860 79520
rect 197640 79410 197650 79480
rect 197850 79410 197860 79480
rect 197640 79360 197860 79410
rect 198140 79590 198360 79640
rect 198140 79520 198150 79590
rect 198350 79520 198360 79590
rect 198140 79480 198360 79520
rect 198140 79410 198150 79480
rect 198350 79410 198360 79480
rect 198140 79360 198360 79410
rect 198640 79590 198860 79640
rect 198640 79520 198650 79590
rect 198850 79520 198860 79590
rect 198640 79480 198860 79520
rect 198640 79410 198650 79480
rect 198850 79410 198860 79480
rect 198640 79360 198860 79410
rect 199140 79590 199360 79640
rect 199140 79520 199150 79590
rect 199350 79520 199360 79590
rect 199140 79480 199360 79520
rect 199140 79410 199150 79480
rect 199350 79410 199360 79480
rect 199140 79360 199360 79410
rect 199640 79590 199860 79640
rect 199640 79520 199650 79590
rect 199850 79520 199860 79590
rect 199640 79480 199860 79520
rect 199640 79410 199650 79480
rect 199850 79410 199860 79480
rect 199640 79360 199860 79410
rect 200140 79590 200360 79640
rect 200140 79520 200150 79590
rect 200350 79520 200360 79590
rect 200140 79480 200360 79520
rect 200140 79410 200150 79480
rect 200350 79410 200360 79480
rect 200140 79360 200360 79410
rect 200640 79590 200860 79640
rect 200640 79520 200650 79590
rect 200850 79520 200860 79590
rect 200640 79480 200860 79520
rect 200640 79410 200650 79480
rect 200850 79410 200860 79480
rect 200640 79360 200860 79410
rect 201140 79590 201360 79640
rect 201140 79520 201150 79590
rect 201350 79520 201360 79590
rect 201140 79480 201360 79520
rect 201140 79410 201150 79480
rect 201350 79410 201360 79480
rect 201140 79360 201360 79410
rect 201640 79590 201860 79640
rect 201640 79520 201650 79590
rect 201850 79520 201860 79590
rect 201640 79480 201860 79520
rect 201640 79410 201650 79480
rect 201850 79410 201860 79480
rect 201640 79360 201860 79410
rect 202140 79590 202360 79640
rect 202140 79520 202150 79590
rect 202350 79520 202360 79590
rect 202140 79480 202360 79520
rect 202140 79410 202150 79480
rect 202350 79410 202360 79480
rect 202140 79360 202360 79410
rect 202640 79590 202860 79640
rect 202640 79520 202650 79590
rect 202850 79520 202860 79590
rect 202640 79480 202860 79520
rect 202640 79410 202650 79480
rect 202850 79410 202860 79480
rect 202640 79360 202860 79410
rect 203140 79590 203360 79640
rect 203140 79520 203150 79590
rect 203350 79520 203360 79590
rect 203140 79480 203360 79520
rect 203140 79410 203150 79480
rect 203350 79410 203360 79480
rect 203140 79360 203360 79410
rect 203640 79590 203860 79640
rect 203640 79520 203650 79590
rect 203850 79520 203860 79590
rect 203640 79480 203860 79520
rect 203640 79410 203650 79480
rect 203850 79410 203860 79480
rect 203640 79360 203860 79410
rect 204140 79590 204360 79640
rect 204140 79520 204150 79590
rect 204350 79520 204360 79590
rect 204140 79480 204360 79520
rect 204140 79410 204150 79480
rect 204350 79410 204360 79480
rect 204140 79360 204360 79410
rect 204640 79590 204860 79640
rect 204640 79520 204650 79590
rect 204850 79520 204860 79590
rect 204640 79480 204860 79520
rect 204640 79410 204650 79480
rect 204850 79410 204860 79480
rect 204640 79360 204860 79410
rect 205140 79590 205360 79640
rect 205140 79520 205150 79590
rect 205350 79520 205360 79590
rect 205140 79480 205360 79520
rect 205140 79410 205150 79480
rect 205350 79410 205360 79480
rect 205140 79360 205360 79410
rect 205640 79590 205860 79640
rect 205640 79520 205650 79590
rect 205850 79520 205860 79590
rect 205640 79480 205860 79520
rect 205640 79410 205650 79480
rect 205850 79410 205860 79480
rect 205640 79360 205860 79410
rect 206140 79590 206360 79640
rect 206140 79520 206150 79590
rect 206350 79520 206360 79590
rect 206140 79480 206360 79520
rect 206140 79410 206150 79480
rect 206350 79410 206360 79480
rect 206140 79360 206360 79410
rect 206640 79590 206860 79640
rect 206640 79520 206650 79590
rect 206850 79520 206860 79590
rect 206640 79480 206860 79520
rect 206640 79410 206650 79480
rect 206850 79410 206860 79480
rect 206640 79360 206860 79410
rect 207140 79590 207360 79640
rect 207140 79520 207150 79590
rect 207350 79520 207360 79590
rect 207140 79480 207360 79520
rect 207140 79410 207150 79480
rect 207350 79410 207360 79480
rect 207140 79360 207360 79410
rect 207640 79590 207860 79640
rect 207640 79520 207650 79590
rect 207850 79520 207860 79590
rect 207640 79480 207860 79520
rect 207640 79410 207650 79480
rect 207850 79410 207860 79480
rect 207640 79360 207860 79410
rect 196000 79350 208000 79360
rect 196000 79150 196020 79350
rect 196090 79150 196410 79350
rect 196480 79150 196520 79350
rect 196590 79150 196910 79350
rect 196980 79150 197020 79350
rect 197090 79150 197410 79350
rect 197480 79150 197520 79350
rect 197590 79150 197910 79350
rect 197980 79150 198020 79350
rect 198090 79150 198410 79350
rect 198480 79150 198520 79350
rect 198590 79150 198910 79350
rect 198980 79150 199020 79350
rect 199090 79150 199410 79350
rect 199480 79150 199520 79350
rect 199590 79150 199910 79350
rect 199980 79150 200020 79350
rect 200090 79150 200410 79350
rect 200480 79150 200520 79350
rect 200590 79150 200910 79350
rect 200980 79150 201020 79350
rect 201090 79150 201410 79350
rect 201480 79150 201520 79350
rect 201590 79150 201910 79350
rect 201980 79150 202020 79350
rect 202090 79150 202410 79350
rect 202480 79150 202520 79350
rect 202590 79150 202910 79350
rect 202980 79150 203020 79350
rect 203090 79150 203410 79350
rect 203480 79150 203520 79350
rect 203590 79150 203910 79350
rect 203980 79150 204020 79350
rect 204090 79150 204410 79350
rect 204480 79150 204520 79350
rect 204590 79150 204910 79350
rect 204980 79150 205020 79350
rect 205090 79150 205410 79350
rect 205480 79150 205520 79350
rect 205590 79150 205910 79350
rect 205980 79150 206020 79350
rect 206090 79150 206410 79350
rect 206480 79150 206520 79350
rect 206590 79150 206910 79350
rect 206980 79150 207020 79350
rect 207090 79150 207410 79350
rect 207480 79150 207520 79350
rect 207590 79150 207910 79350
rect 207980 79150 208000 79350
rect 196000 79140 208000 79150
rect 196140 79090 196360 79140
rect 196140 79020 196150 79090
rect 196350 79020 196360 79090
rect 196140 78980 196360 79020
rect 196140 78910 196150 78980
rect 196350 78910 196360 78980
rect 196140 78860 196360 78910
rect 196640 79090 196860 79140
rect 196640 79020 196650 79090
rect 196850 79020 196860 79090
rect 196640 78980 196860 79020
rect 196640 78910 196650 78980
rect 196850 78910 196860 78980
rect 196640 78860 196860 78910
rect 197140 79090 197360 79140
rect 197140 79020 197150 79090
rect 197350 79020 197360 79090
rect 197140 78980 197360 79020
rect 197140 78910 197150 78980
rect 197350 78910 197360 78980
rect 197140 78860 197360 78910
rect 197640 79090 197860 79140
rect 197640 79020 197650 79090
rect 197850 79020 197860 79090
rect 197640 78980 197860 79020
rect 197640 78910 197650 78980
rect 197850 78910 197860 78980
rect 197640 78860 197860 78910
rect 198140 79090 198360 79140
rect 198140 79020 198150 79090
rect 198350 79020 198360 79090
rect 198140 78980 198360 79020
rect 198140 78910 198150 78980
rect 198350 78910 198360 78980
rect 198140 78860 198360 78910
rect 198640 79090 198860 79140
rect 198640 79020 198650 79090
rect 198850 79020 198860 79090
rect 198640 78980 198860 79020
rect 198640 78910 198650 78980
rect 198850 78910 198860 78980
rect 198640 78860 198860 78910
rect 199140 79090 199360 79140
rect 199140 79020 199150 79090
rect 199350 79020 199360 79090
rect 199140 78980 199360 79020
rect 199140 78910 199150 78980
rect 199350 78910 199360 78980
rect 199140 78860 199360 78910
rect 199640 79090 199860 79140
rect 199640 79020 199650 79090
rect 199850 79020 199860 79090
rect 199640 78980 199860 79020
rect 199640 78910 199650 78980
rect 199850 78910 199860 78980
rect 199640 78860 199860 78910
rect 200140 79090 200360 79140
rect 200140 79020 200150 79090
rect 200350 79020 200360 79090
rect 200140 78980 200360 79020
rect 200140 78910 200150 78980
rect 200350 78910 200360 78980
rect 200140 78860 200360 78910
rect 200640 79090 200860 79140
rect 200640 79020 200650 79090
rect 200850 79020 200860 79090
rect 200640 78980 200860 79020
rect 200640 78910 200650 78980
rect 200850 78910 200860 78980
rect 200640 78860 200860 78910
rect 201140 79090 201360 79140
rect 201140 79020 201150 79090
rect 201350 79020 201360 79090
rect 201140 78980 201360 79020
rect 201140 78910 201150 78980
rect 201350 78910 201360 78980
rect 201140 78860 201360 78910
rect 201640 79090 201860 79140
rect 201640 79020 201650 79090
rect 201850 79020 201860 79090
rect 201640 78980 201860 79020
rect 201640 78910 201650 78980
rect 201850 78910 201860 78980
rect 201640 78860 201860 78910
rect 202140 79090 202360 79140
rect 202140 79020 202150 79090
rect 202350 79020 202360 79090
rect 202140 78980 202360 79020
rect 202140 78910 202150 78980
rect 202350 78910 202360 78980
rect 202140 78860 202360 78910
rect 202640 79090 202860 79140
rect 202640 79020 202650 79090
rect 202850 79020 202860 79090
rect 202640 78980 202860 79020
rect 202640 78910 202650 78980
rect 202850 78910 202860 78980
rect 202640 78860 202860 78910
rect 203140 79090 203360 79140
rect 203140 79020 203150 79090
rect 203350 79020 203360 79090
rect 203140 78980 203360 79020
rect 203140 78910 203150 78980
rect 203350 78910 203360 78980
rect 203140 78860 203360 78910
rect 203640 79090 203860 79140
rect 203640 79020 203650 79090
rect 203850 79020 203860 79090
rect 203640 78980 203860 79020
rect 203640 78910 203650 78980
rect 203850 78910 203860 78980
rect 203640 78860 203860 78910
rect 204140 79090 204360 79140
rect 204140 79020 204150 79090
rect 204350 79020 204360 79090
rect 204140 78980 204360 79020
rect 204140 78910 204150 78980
rect 204350 78910 204360 78980
rect 204140 78860 204360 78910
rect 204640 79090 204860 79140
rect 204640 79020 204650 79090
rect 204850 79020 204860 79090
rect 204640 78980 204860 79020
rect 204640 78910 204650 78980
rect 204850 78910 204860 78980
rect 204640 78860 204860 78910
rect 205140 79090 205360 79140
rect 205140 79020 205150 79090
rect 205350 79020 205360 79090
rect 205140 78980 205360 79020
rect 205140 78910 205150 78980
rect 205350 78910 205360 78980
rect 205140 78860 205360 78910
rect 205640 79090 205860 79140
rect 205640 79020 205650 79090
rect 205850 79020 205860 79090
rect 205640 78980 205860 79020
rect 205640 78910 205650 78980
rect 205850 78910 205860 78980
rect 205640 78860 205860 78910
rect 206140 79090 206360 79140
rect 206140 79020 206150 79090
rect 206350 79020 206360 79090
rect 206140 78980 206360 79020
rect 206140 78910 206150 78980
rect 206350 78910 206360 78980
rect 206140 78860 206360 78910
rect 206640 79090 206860 79140
rect 206640 79020 206650 79090
rect 206850 79020 206860 79090
rect 206640 78980 206860 79020
rect 206640 78910 206650 78980
rect 206850 78910 206860 78980
rect 206640 78860 206860 78910
rect 207140 79090 207360 79140
rect 207140 79020 207150 79090
rect 207350 79020 207360 79090
rect 207140 78980 207360 79020
rect 207140 78910 207150 78980
rect 207350 78910 207360 78980
rect 207140 78860 207360 78910
rect 207640 79090 207860 79140
rect 207640 79020 207650 79090
rect 207850 79020 207860 79090
rect 207640 78980 207860 79020
rect 207640 78910 207650 78980
rect 207850 78910 207860 78980
rect 207640 78860 207860 78910
rect 196000 78850 208000 78860
rect 196000 78650 196020 78850
rect 196090 78650 196410 78850
rect 196480 78650 196520 78850
rect 196590 78650 196910 78850
rect 196980 78650 197020 78850
rect 197090 78650 197410 78850
rect 197480 78650 197520 78850
rect 197590 78650 197910 78850
rect 197980 78650 198020 78850
rect 198090 78650 198410 78850
rect 198480 78650 198520 78850
rect 198590 78650 198910 78850
rect 198980 78650 199020 78850
rect 199090 78650 199410 78850
rect 199480 78650 199520 78850
rect 199590 78650 199910 78850
rect 199980 78650 200020 78850
rect 200090 78650 200410 78850
rect 200480 78650 200520 78850
rect 200590 78650 200910 78850
rect 200980 78650 201020 78850
rect 201090 78650 201410 78850
rect 201480 78650 201520 78850
rect 201590 78650 201910 78850
rect 201980 78650 202020 78850
rect 202090 78650 202410 78850
rect 202480 78650 202520 78850
rect 202590 78650 202910 78850
rect 202980 78650 203020 78850
rect 203090 78650 203410 78850
rect 203480 78650 203520 78850
rect 203590 78650 203910 78850
rect 203980 78650 204020 78850
rect 204090 78650 204410 78850
rect 204480 78650 204520 78850
rect 204590 78650 204910 78850
rect 204980 78650 205020 78850
rect 205090 78650 205410 78850
rect 205480 78650 205520 78850
rect 205590 78650 205910 78850
rect 205980 78650 206020 78850
rect 206090 78650 206410 78850
rect 206480 78650 206520 78850
rect 206590 78650 206910 78850
rect 206980 78650 207020 78850
rect 207090 78650 207410 78850
rect 207480 78650 207520 78850
rect 207590 78650 207910 78850
rect 207980 78650 208000 78850
rect 196000 78640 208000 78650
rect 196140 78590 196360 78640
rect 196140 78520 196150 78590
rect 196350 78520 196360 78590
rect 196140 78480 196360 78520
rect 196140 78410 196150 78480
rect 196350 78410 196360 78480
rect 196140 78360 196360 78410
rect 196640 78590 196860 78640
rect 196640 78520 196650 78590
rect 196850 78520 196860 78590
rect 196640 78480 196860 78520
rect 196640 78410 196650 78480
rect 196850 78410 196860 78480
rect 196640 78360 196860 78410
rect 197140 78590 197360 78640
rect 197140 78520 197150 78590
rect 197350 78520 197360 78590
rect 197140 78480 197360 78520
rect 197140 78410 197150 78480
rect 197350 78410 197360 78480
rect 197140 78360 197360 78410
rect 197640 78590 197860 78640
rect 197640 78520 197650 78590
rect 197850 78520 197860 78590
rect 197640 78480 197860 78520
rect 197640 78410 197650 78480
rect 197850 78410 197860 78480
rect 197640 78360 197860 78410
rect 198140 78590 198360 78640
rect 198140 78520 198150 78590
rect 198350 78520 198360 78590
rect 198140 78480 198360 78520
rect 198140 78410 198150 78480
rect 198350 78410 198360 78480
rect 198140 78360 198360 78410
rect 198640 78590 198860 78640
rect 198640 78520 198650 78590
rect 198850 78520 198860 78590
rect 198640 78480 198860 78520
rect 198640 78410 198650 78480
rect 198850 78410 198860 78480
rect 198640 78360 198860 78410
rect 199140 78590 199360 78640
rect 199140 78520 199150 78590
rect 199350 78520 199360 78590
rect 199140 78480 199360 78520
rect 199140 78410 199150 78480
rect 199350 78410 199360 78480
rect 199140 78360 199360 78410
rect 199640 78590 199860 78640
rect 199640 78520 199650 78590
rect 199850 78520 199860 78590
rect 199640 78480 199860 78520
rect 199640 78410 199650 78480
rect 199850 78410 199860 78480
rect 199640 78360 199860 78410
rect 200140 78590 200360 78640
rect 200140 78520 200150 78590
rect 200350 78520 200360 78590
rect 200140 78480 200360 78520
rect 200140 78410 200150 78480
rect 200350 78410 200360 78480
rect 200140 78360 200360 78410
rect 200640 78590 200860 78640
rect 200640 78520 200650 78590
rect 200850 78520 200860 78590
rect 200640 78480 200860 78520
rect 200640 78410 200650 78480
rect 200850 78410 200860 78480
rect 200640 78360 200860 78410
rect 201140 78590 201360 78640
rect 201140 78520 201150 78590
rect 201350 78520 201360 78590
rect 201140 78480 201360 78520
rect 201140 78410 201150 78480
rect 201350 78410 201360 78480
rect 201140 78360 201360 78410
rect 201640 78590 201860 78640
rect 201640 78520 201650 78590
rect 201850 78520 201860 78590
rect 201640 78480 201860 78520
rect 201640 78410 201650 78480
rect 201850 78410 201860 78480
rect 201640 78360 201860 78410
rect 202140 78590 202360 78640
rect 202140 78520 202150 78590
rect 202350 78520 202360 78590
rect 202140 78480 202360 78520
rect 202140 78410 202150 78480
rect 202350 78410 202360 78480
rect 202140 78360 202360 78410
rect 202640 78590 202860 78640
rect 202640 78520 202650 78590
rect 202850 78520 202860 78590
rect 202640 78480 202860 78520
rect 202640 78410 202650 78480
rect 202850 78410 202860 78480
rect 202640 78360 202860 78410
rect 203140 78590 203360 78640
rect 203140 78520 203150 78590
rect 203350 78520 203360 78590
rect 203140 78480 203360 78520
rect 203140 78410 203150 78480
rect 203350 78410 203360 78480
rect 203140 78360 203360 78410
rect 203640 78590 203860 78640
rect 203640 78520 203650 78590
rect 203850 78520 203860 78590
rect 203640 78480 203860 78520
rect 203640 78410 203650 78480
rect 203850 78410 203860 78480
rect 203640 78360 203860 78410
rect 204140 78590 204360 78640
rect 204140 78520 204150 78590
rect 204350 78520 204360 78590
rect 204140 78480 204360 78520
rect 204140 78410 204150 78480
rect 204350 78410 204360 78480
rect 204140 78360 204360 78410
rect 204640 78590 204860 78640
rect 204640 78520 204650 78590
rect 204850 78520 204860 78590
rect 204640 78480 204860 78520
rect 204640 78410 204650 78480
rect 204850 78410 204860 78480
rect 204640 78360 204860 78410
rect 205140 78590 205360 78640
rect 205140 78520 205150 78590
rect 205350 78520 205360 78590
rect 205140 78480 205360 78520
rect 205140 78410 205150 78480
rect 205350 78410 205360 78480
rect 205140 78360 205360 78410
rect 205640 78590 205860 78640
rect 205640 78520 205650 78590
rect 205850 78520 205860 78590
rect 205640 78480 205860 78520
rect 205640 78410 205650 78480
rect 205850 78410 205860 78480
rect 205640 78360 205860 78410
rect 206140 78590 206360 78640
rect 206140 78520 206150 78590
rect 206350 78520 206360 78590
rect 206140 78480 206360 78520
rect 206140 78410 206150 78480
rect 206350 78410 206360 78480
rect 206140 78360 206360 78410
rect 206640 78590 206860 78640
rect 206640 78520 206650 78590
rect 206850 78520 206860 78590
rect 206640 78480 206860 78520
rect 206640 78410 206650 78480
rect 206850 78410 206860 78480
rect 206640 78360 206860 78410
rect 207140 78590 207360 78640
rect 207140 78520 207150 78590
rect 207350 78520 207360 78590
rect 207140 78480 207360 78520
rect 207140 78410 207150 78480
rect 207350 78410 207360 78480
rect 207140 78360 207360 78410
rect 207640 78590 207860 78640
rect 207640 78520 207650 78590
rect 207850 78520 207860 78590
rect 207640 78480 207860 78520
rect 207640 78410 207650 78480
rect 207850 78410 207860 78480
rect 207640 78360 207860 78410
rect 196000 78350 208000 78360
rect 196000 78150 196020 78350
rect 196090 78150 196410 78350
rect 196480 78150 196520 78350
rect 196590 78150 196910 78350
rect 196980 78150 197020 78350
rect 197090 78150 197410 78350
rect 197480 78150 197520 78350
rect 197590 78150 197910 78350
rect 197980 78150 198020 78350
rect 198090 78150 198410 78350
rect 198480 78150 198520 78350
rect 198590 78150 198910 78350
rect 198980 78150 199020 78350
rect 199090 78150 199410 78350
rect 199480 78150 199520 78350
rect 199590 78150 199910 78350
rect 199980 78150 200020 78350
rect 200090 78150 200410 78350
rect 200480 78150 200520 78350
rect 200590 78150 200910 78350
rect 200980 78150 201020 78350
rect 201090 78150 201410 78350
rect 201480 78150 201520 78350
rect 201590 78150 201910 78350
rect 201980 78150 202020 78350
rect 202090 78150 202410 78350
rect 202480 78150 202520 78350
rect 202590 78150 202910 78350
rect 202980 78150 203020 78350
rect 203090 78150 203410 78350
rect 203480 78150 203520 78350
rect 203590 78150 203910 78350
rect 203980 78150 204020 78350
rect 204090 78150 204410 78350
rect 204480 78150 204520 78350
rect 204590 78150 204910 78350
rect 204980 78150 205020 78350
rect 205090 78150 205410 78350
rect 205480 78150 205520 78350
rect 205590 78150 205910 78350
rect 205980 78150 206020 78350
rect 206090 78150 206410 78350
rect 206480 78150 206520 78350
rect 206590 78150 206910 78350
rect 206980 78150 207020 78350
rect 207090 78150 207410 78350
rect 207480 78150 207520 78350
rect 207590 78150 207910 78350
rect 207980 78150 208000 78350
rect 196000 78140 208000 78150
rect 196140 78090 196360 78140
rect 196140 78020 196150 78090
rect 196350 78020 196360 78090
rect 196140 77980 196360 78020
rect 196140 77910 196150 77980
rect 196350 77910 196360 77980
rect 196140 77860 196360 77910
rect 196640 78090 196860 78140
rect 196640 78020 196650 78090
rect 196850 78020 196860 78090
rect 196640 77980 196860 78020
rect 196640 77910 196650 77980
rect 196850 77910 196860 77980
rect 196640 77860 196860 77910
rect 197140 78090 197360 78140
rect 197140 78020 197150 78090
rect 197350 78020 197360 78090
rect 197140 77980 197360 78020
rect 197140 77910 197150 77980
rect 197350 77910 197360 77980
rect 197140 77860 197360 77910
rect 197640 78090 197860 78140
rect 197640 78020 197650 78090
rect 197850 78020 197860 78090
rect 197640 77980 197860 78020
rect 197640 77910 197650 77980
rect 197850 77910 197860 77980
rect 197640 77860 197860 77910
rect 198140 78090 198360 78140
rect 198140 78020 198150 78090
rect 198350 78020 198360 78090
rect 198140 77980 198360 78020
rect 198140 77910 198150 77980
rect 198350 77910 198360 77980
rect 198140 77860 198360 77910
rect 198640 78090 198860 78140
rect 198640 78020 198650 78090
rect 198850 78020 198860 78090
rect 198640 77980 198860 78020
rect 198640 77910 198650 77980
rect 198850 77910 198860 77980
rect 198640 77860 198860 77910
rect 199140 78090 199360 78140
rect 199140 78020 199150 78090
rect 199350 78020 199360 78090
rect 199140 77980 199360 78020
rect 199140 77910 199150 77980
rect 199350 77910 199360 77980
rect 199140 77860 199360 77910
rect 199640 78090 199860 78140
rect 199640 78020 199650 78090
rect 199850 78020 199860 78090
rect 199640 77980 199860 78020
rect 199640 77910 199650 77980
rect 199850 77910 199860 77980
rect 199640 77860 199860 77910
rect 200140 78090 200360 78140
rect 200140 78020 200150 78090
rect 200350 78020 200360 78090
rect 200140 77980 200360 78020
rect 200140 77910 200150 77980
rect 200350 77910 200360 77980
rect 200140 77860 200360 77910
rect 200640 78090 200860 78140
rect 200640 78020 200650 78090
rect 200850 78020 200860 78090
rect 200640 77980 200860 78020
rect 200640 77910 200650 77980
rect 200850 77910 200860 77980
rect 200640 77860 200860 77910
rect 201140 78090 201360 78140
rect 201140 78020 201150 78090
rect 201350 78020 201360 78090
rect 201140 77980 201360 78020
rect 201140 77910 201150 77980
rect 201350 77910 201360 77980
rect 201140 77860 201360 77910
rect 201640 78090 201860 78140
rect 201640 78020 201650 78090
rect 201850 78020 201860 78090
rect 201640 77980 201860 78020
rect 201640 77910 201650 77980
rect 201850 77910 201860 77980
rect 201640 77860 201860 77910
rect 202140 78090 202360 78140
rect 202140 78020 202150 78090
rect 202350 78020 202360 78090
rect 202140 77980 202360 78020
rect 202140 77910 202150 77980
rect 202350 77910 202360 77980
rect 202140 77860 202360 77910
rect 202640 78090 202860 78140
rect 202640 78020 202650 78090
rect 202850 78020 202860 78090
rect 202640 77980 202860 78020
rect 202640 77910 202650 77980
rect 202850 77910 202860 77980
rect 202640 77860 202860 77910
rect 203140 78090 203360 78140
rect 203140 78020 203150 78090
rect 203350 78020 203360 78090
rect 203140 77980 203360 78020
rect 203140 77910 203150 77980
rect 203350 77910 203360 77980
rect 203140 77860 203360 77910
rect 203640 78090 203860 78140
rect 203640 78020 203650 78090
rect 203850 78020 203860 78090
rect 203640 77980 203860 78020
rect 203640 77910 203650 77980
rect 203850 77910 203860 77980
rect 203640 77860 203860 77910
rect 204140 78090 204360 78140
rect 204140 78020 204150 78090
rect 204350 78020 204360 78090
rect 204140 77980 204360 78020
rect 204140 77910 204150 77980
rect 204350 77910 204360 77980
rect 204140 77860 204360 77910
rect 204640 78090 204860 78140
rect 204640 78020 204650 78090
rect 204850 78020 204860 78090
rect 204640 77980 204860 78020
rect 204640 77910 204650 77980
rect 204850 77910 204860 77980
rect 204640 77860 204860 77910
rect 205140 78090 205360 78140
rect 205140 78020 205150 78090
rect 205350 78020 205360 78090
rect 205140 77980 205360 78020
rect 205140 77910 205150 77980
rect 205350 77910 205360 77980
rect 205140 77860 205360 77910
rect 205640 78090 205860 78140
rect 205640 78020 205650 78090
rect 205850 78020 205860 78090
rect 205640 77980 205860 78020
rect 205640 77910 205650 77980
rect 205850 77910 205860 77980
rect 205640 77860 205860 77910
rect 206140 78090 206360 78140
rect 206140 78020 206150 78090
rect 206350 78020 206360 78090
rect 206140 77980 206360 78020
rect 206140 77910 206150 77980
rect 206350 77910 206360 77980
rect 206140 77860 206360 77910
rect 206640 78090 206860 78140
rect 206640 78020 206650 78090
rect 206850 78020 206860 78090
rect 206640 77980 206860 78020
rect 206640 77910 206650 77980
rect 206850 77910 206860 77980
rect 206640 77860 206860 77910
rect 207140 78090 207360 78140
rect 207140 78020 207150 78090
rect 207350 78020 207360 78090
rect 207140 77980 207360 78020
rect 207140 77910 207150 77980
rect 207350 77910 207360 77980
rect 207140 77860 207360 77910
rect 207640 78090 207860 78140
rect 207640 78020 207650 78090
rect 207850 78020 207860 78090
rect 207640 77980 207860 78020
rect 207640 77910 207650 77980
rect 207850 77910 207860 77980
rect 207640 77860 207860 77910
rect 196000 77850 208000 77860
rect 196000 77650 196020 77850
rect 196090 77650 196410 77850
rect 196480 77650 196520 77850
rect 196590 77650 196910 77850
rect 196980 77650 197020 77850
rect 197090 77650 197410 77850
rect 197480 77650 197520 77850
rect 197590 77650 197910 77850
rect 197980 77650 198020 77850
rect 198090 77650 198410 77850
rect 198480 77650 198520 77850
rect 198590 77650 198910 77850
rect 198980 77650 199020 77850
rect 199090 77650 199410 77850
rect 199480 77650 199520 77850
rect 199590 77650 199910 77850
rect 199980 77650 200020 77850
rect 200090 77650 200410 77850
rect 200480 77650 200520 77850
rect 200590 77650 200910 77850
rect 200980 77650 201020 77850
rect 201090 77650 201410 77850
rect 201480 77650 201520 77850
rect 201590 77650 201910 77850
rect 201980 77650 202020 77850
rect 202090 77650 202410 77850
rect 202480 77650 202520 77850
rect 202590 77650 202910 77850
rect 202980 77650 203020 77850
rect 203090 77650 203410 77850
rect 203480 77650 203520 77850
rect 203590 77650 203910 77850
rect 203980 77650 204020 77850
rect 204090 77650 204410 77850
rect 204480 77650 204520 77850
rect 204590 77650 204910 77850
rect 204980 77650 205020 77850
rect 205090 77650 205410 77850
rect 205480 77650 205520 77850
rect 205590 77650 205910 77850
rect 205980 77650 206020 77850
rect 206090 77650 206410 77850
rect 206480 77650 206520 77850
rect 206590 77650 206910 77850
rect 206980 77650 207020 77850
rect 207090 77650 207410 77850
rect 207480 77650 207520 77850
rect 207590 77650 207910 77850
rect 207980 77650 208000 77850
rect 196000 77640 208000 77650
rect 196140 77590 196360 77640
rect 196140 77520 196150 77590
rect 196350 77520 196360 77590
rect 196140 77480 196360 77520
rect 196140 77410 196150 77480
rect 196350 77410 196360 77480
rect 196140 77360 196360 77410
rect 196640 77590 196860 77640
rect 196640 77520 196650 77590
rect 196850 77520 196860 77590
rect 196640 77480 196860 77520
rect 196640 77410 196650 77480
rect 196850 77410 196860 77480
rect 196640 77360 196860 77410
rect 197140 77590 197360 77640
rect 197140 77520 197150 77590
rect 197350 77520 197360 77590
rect 197140 77480 197360 77520
rect 197140 77410 197150 77480
rect 197350 77410 197360 77480
rect 197140 77360 197360 77410
rect 197640 77590 197860 77640
rect 197640 77520 197650 77590
rect 197850 77520 197860 77590
rect 197640 77480 197860 77520
rect 197640 77410 197650 77480
rect 197850 77410 197860 77480
rect 197640 77360 197860 77410
rect 198140 77590 198360 77640
rect 198140 77520 198150 77590
rect 198350 77520 198360 77590
rect 198140 77480 198360 77520
rect 198140 77410 198150 77480
rect 198350 77410 198360 77480
rect 198140 77360 198360 77410
rect 198640 77590 198860 77640
rect 198640 77520 198650 77590
rect 198850 77520 198860 77590
rect 198640 77480 198860 77520
rect 198640 77410 198650 77480
rect 198850 77410 198860 77480
rect 198640 77360 198860 77410
rect 199140 77590 199360 77640
rect 199140 77520 199150 77590
rect 199350 77520 199360 77590
rect 199140 77480 199360 77520
rect 199140 77410 199150 77480
rect 199350 77410 199360 77480
rect 199140 77360 199360 77410
rect 199640 77590 199860 77640
rect 199640 77520 199650 77590
rect 199850 77520 199860 77590
rect 199640 77480 199860 77520
rect 199640 77410 199650 77480
rect 199850 77410 199860 77480
rect 199640 77360 199860 77410
rect 200140 77590 200360 77640
rect 200140 77520 200150 77590
rect 200350 77520 200360 77590
rect 200140 77480 200360 77520
rect 200140 77410 200150 77480
rect 200350 77410 200360 77480
rect 200140 77360 200360 77410
rect 200640 77590 200860 77640
rect 200640 77520 200650 77590
rect 200850 77520 200860 77590
rect 200640 77480 200860 77520
rect 200640 77410 200650 77480
rect 200850 77410 200860 77480
rect 200640 77360 200860 77410
rect 201140 77590 201360 77640
rect 201140 77520 201150 77590
rect 201350 77520 201360 77590
rect 201140 77480 201360 77520
rect 201140 77410 201150 77480
rect 201350 77410 201360 77480
rect 201140 77360 201360 77410
rect 201640 77590 201860 77640
rect 201640 77520 201650 77590
rect 201850 77520 201860 77590
rect 201640 77480 201860 77520
rect 201640 77410 201650 77480
rect 201850 77410 201860 77480
rect 201640 77360 201860 77410
rect 202140 77590 202360 77640
rect 202140 77520 202150 77590
rect 202350 77520 202360 77590
rect 202140 77480 202360 77520
rect 202140 77410 202150 77480
rect 202350 77410 202360 77480
rect 202140 77360 202360 77410
rect 202640 77590 202860 77640
rect 202640 77520 202650 77590
rect 202850 77520 202860 77590
rect 202640 77480 202860 77520
rect 202640 77410 202650 77480
rect 202850 77410 202860 77480
rect 202640 77360 202860 77410
rect 203140 77590 203360 77640
rect 203140 77520 203150 77590
rect 203350 77520 203360 77590
rect 203140 77480 203360 77520
rect 203140 77410 203150 77480
rect 203350 77410 203360 77480
rect 203140 77360 203360 77410
rect 203640 77590 203860 77640
rect 203640 77520 203650 77590
rect 203850 77520 203860 77590
rect 203640 77480 203860 77520
rect 203640 77410 203650 77480
rect 203850 77410 203860 77480
rect 203640 77360 203860 77410
rect 204140 77590 204360 77640
rect 204140 77520 204150 77590
rect 204350 77520 204360 77590
rect 204140 77480 204360 77520
rect 204140 77410 204150 77480
rect 204350 77410 204360 77480
rect 204140 77360 204360 77410
rect 204640 77590 204860 77640
rect 204640 77520 204650 77590
rect 204850 77520 204860 77590
rect 204640 77480 204860 77520
rect 204640 77410 204650 77480
rect 204850 77410 204860 77480
rect 204640 77360 204860 77410
rect 205140 77590 205360 77640
rect 205140 77520 205150 77590
rect 205350 77520 205360 77590
rect 205140 77480 205360 77520
rect 205140 77410 205150 77480
rect 205350 77410 205360 77480
rect 205140 77360 205360 77410
rect 205640 77590 205860 77640
rect 205640 77520 205650 77590
rect 205850 77520 205860 77590
rect 205640 77480 205860 77520
rect 205640 77410 205650 77480
rect 205850 77410 205860 77480
rect 205640 77360 205860 77410
rect 206140 77590 206360 77640
rect 206140 77520 206150 77590
rect 206350 77520 206360 77590
rect 206140 77480 206360 77520
rect 206140 77410 206150 77480
rect 206350 77410 206360 77480
rect 206140 77360 206360 77410
rect 206640 77590 206860 77640
rect 206640 77520 206650 77590
rect 206850 77520 206860 77590
rect 206640 77480 206860 77520
rect 206640 77410 206650 77480
rect 206850 77410 206860 77480
rect 206640 77360 206860 77410
rect 207140 77590 207360 77640
rect 207140 77520 207150 77590
rect 207350 77520 207360 77590
rect 207140 77480 207360 77520
rect 207140 77410 207150 77480
rect 207350 77410 207360 77480
rect 207140 77360 207360 77410
rect 207640 77590 207860 77640
rect 207640 77520 207650 77590
rect 207850 77520 207860 77590
rect 207640 77480 207860 77520
rect 207640 77410 207650 77480
rect 207850 77410 207860 77480
rect 207640 77360 207860 77410
rect 196000 77350 208000 77360
rect 196000 77150 196020 77350
rect 196090 77150 196410 77350
rect 196480 77150 196520 77350
rect 196590 77150 196910 77350
rect 196980 77150 197020 77350
rect 197090 77150 197410 77350
rect 197480 77150 197520 77350
rect 197590 77150 197910 77350
rect 197980 77150 198020 77350
rect 198090 77150 198410 77350
rect 198480 77150 198520 77350
rect 198590 77150 198910 77350
rect 198980 77150 199020 77350
rect 199090 77150 199410 77350
rect 199480 77150 199520 77350
rect 199590 77150 199910 77350
rect 199980 77150 200020 77350
rect 200090 77150 200410 77350
rect 200480 77150 200520 77350
rect 200590 77150 200910 77350
rect 200980 77150 201020 77350
rect 201090 77150 201410 77350
rect 201480 77150 201520 77350
rect 201590 77150 201910 77350
rect 201980 77150 202020 77350
rect 202090 77150 202410 77350
rect 202480 77150 202520 77350
rect 202590 77150 202910 77350
rect 202980 77150 203020 77350
rect 203090 77150 203410 77350
rect 203480 77150 203520 77350
rect 203590 77150 203910 77350
rect 203980 77150 204020 77350
rect 204090 77150 204410 77350
rect 204480 77150 204520 77350
rect 204590 77150 204910 77350
rect 204980 77150 205020 77350
rect 205090 77150 205410 77350
rect 205480 77150 205520 77350
rect 205590 77150 205910 77350
rect 205980 77150 206020 77350
rect 206090 77150 206410 77350
rect 206480 77150 206520 77350
rect 206590 77150 206910 77350
rect 206980 77150 207020 77350
rect 207090 77150 207410 77350
rect 207480 77150 207520 77350
rect 207590 77150 207910 77350
rect 207980 77150 208000 77350
rect 196000 77140 208000 77150
rect 196140 77090 196360 77140
rect 196140 77020 196150 77090
rect 196350 77020 196360 77090
rect 196140 76980 196360 77020
rect 196140 76910 196150 76980
rect 196350 76910 196360 76980
rect 196140 76860 196360 76910
rect 196640 77090 196860 77140
rect 196640 77020 196650 77090
rect 196850 77020 196860 77090
rect 196640 76980 196860 77020
rect 196640 76910 196650 76980
rect 196850 76910 196860 76980
rect 196640 76860 196860 76910
rect 197140 77090 197360 77140
rect 197140 77020 197150 77090
rect 197350 77020 197360 77090
rect 197140 76980 197360 77020
rect 197140 76910 197150 76980
rect 197350 76910 197360 76980
rect 197140 76860 197360 76910
rect 197640 77090 197860 77140
rect 197640 77020 197650 77090
rect 197850 77020 197860 77090
rect 197640 76980 197860 77020
rect 197640 76910 197650 76980
rect 197850 76910 197860 76980
rect 197640 76860 197860 76910
rect 198140 77090 198360 77140
rect 198140 77020 198150 77090
rect 198350 77020 198360 77090
rect 198140 76980 198360 77020
rect 198140 76910 198150 76980
rect 198350 76910 198360 76980
rect 198140 76860 198360 76910
rect 198640 77090 198860 77140
rect 198640 77020 198650 77090
rect 198850 77020 198860 77090
rect 198640 76980 198860 77020
rect 198640 76910 198650 76980
rect 198850 76910 198860 76980
rect 198640 76860 198860 76910
rect 199140 77090 199360 77140
rect 199140 77020 199150 77090
rect 199350 77020 199360 77090
rect 199140 76980 199360 77020
rect 199140 76910 199150 76980
rect 199350 76910 199360 76980
rect 199140 76860 199360 76910
rect 199640 77090 199860 77140
rect 199640 77020 199650 77090
rect 199850 77020 199860 77090
rect 199640 76980 199860 77020
rect 199640 76910 199650 76980
rect 199850 76910 199860 76980
rect 199640 76860 199860 76910
rect 200140 77090 200360 77140
rect 200140 77020 200150 77090
rect 200350 77020 200360 77090
rect 200140 76980 200360 77020
rect 200140 76910 200150 76980
rect 200350 76910 200360 76980
rect 200140 76860 200360 76910
rect 200640 77090 200860 77140
rect 200640 77020 200650 77090
rect 200850 77020 200860 77090
rect 200640 76980 200860 77020
rect 200640 76910 200650 76980
rect 200850 76910 200860 76980
rect 200640 76860 200860 76910
rect 201140 77090 201360 77140
rect 201140 77020 201150 77090
rect 201350 77020 201360 77090
rect 201140 76980 201360 77020
rect 201140 76910 201150 76980
rect 201350 76910 201360 76980
rect 201140 76860 201360 76910
rect 201640 77090 201860 77140
rect 201640 77020 201650 77090
rect 201850 77020 201860 77090
rect 201640 76980 201860 77020
rect 201640 76910 201650 76980
rect 201850 76910 201860 76980
rect 201640 76860 201860 76910
rect 202140 77090 202360 77140
rect 202140 77020 202150 77090
rect 202350 77020 202360 77090
rect 202140 76980 202360 77020
rect 202140 76910 202150 76980
rect 202350 76910 202360 76980
rect 202140 76860 202360 76910
rect 202640 77090 202860 77140
rect 202640 77020 202650 77090
rect 202850 77020 202860 77090
rect 202640 76980 202860 77020
rect 202640 76910 202650 76980
rect 202850 76910 202860 76980
rect 202640 76860 202860 76910
rect 203140 77090 203360 77140
rect 203140 77020 203150 77090
rect 203350 77020 203360 77090
rect 203140 76980 203360 77020
rect 203140 76910 203150 76980
rect 203350 76910 203360 76980
rect 203140 76860 203360 76910
rect 203640 77090 203860 77140
rect 203640 77020 203650 77090
rect 203850 77020 203860 77090
rect 203640 76980 203860 77020
rect 203640 76910 203650 76980
rect 203850 76910 203860 76980
rect 203640 76860 203860 76910
rect 204140 77090 204360 77140
rect 204140 77020 204150 77090
rect 204350 77020 204360 77090
rect 204140 76980 204360 77020
rect 204140 76910 204150 76980
rect 204350 76910 204360 76980
rect 204140 76860 204360 76910
rect 204640 77090 204860 77140
rect 204640 77020 204650 77090
rect 204850 77020 204860 77090
rect 204640 76980 204860 77020
rect 204640 76910 204650 76980
rect 204850 76910 204860 76980
rect 204640 76860 204860 76910
rect 205140 77090 205360 77140
rect 205140 77020 205150 77090
rect 205350 77020 205360 77090
rect 205140 76980 205360 77020
rect 205140 76910 205150 76980
rect 205350 76910 205360 76980
rect 205140 76860 205360 76910
rect 205640 77090 205860 77140
rect 205640 77020 205650 77090
rect 205850 77020 205860 77090
rect 205640 76980 205860 77020
rect 205640 76910 205650 76980
rect 205850 76910 205860 76980
rect 205640 76860 205860 76910
rect 206140 77090 206360 77140
rect 206140 77020 206150 77090
rect 206350 77020 206360 77090
rect 206140 76980 206360 77020
rect 206140 76910 206150 76980
rect 206350 76910 206360 76980
rect 206140 76860 206360 76910
rect 206640 77090 206860 77140
rect 206640 77020 206650 77090
rect 206850 77020 206860 77090
rect 206640 76980 206860 77020
rect 206640 76910 206650 76980
rect 206850 76910 206860 76980
rect 206640 76860 206860 76910
rect 207140 77090 207360 77140
rect 207140 77020 207150 77090
rect 207350 77020 207360 77090
rect 207140 76980 207360 77020
rect 207140 76910 207150 76980
rect 207350 76910 207360 76980
rect 207140 76860 207360 76910
rect 207640 77090 207860 77140
rect 207640 77020 207650 77090
rect 207850 77020 207860 77090
rect 207640 76980 207860 77020
rect 207640 76910 207650 76980
rect 207850 76910 207860 76980
rect 207640 76860 207860 76910
rect 196000 76850 208000 76860
rect 196000 76650 196020 76850
rect 196090 76650 196410 76850
rect 196480 76650 196520 76850
rect 196590 76650 196910 76850
rect 196980 76650 197020 76850
rect 197090 76650 197410 76850
rect 197480 76650 197520 76850
rect 197590 76650 197910 76850
rect 197980 76650 198020 76850
rect 198090 76650 198410 76850
rect 198480 76650 198520 76850
rect 198590 76650 198910 76850
rect 198980 76650 199020 76850
rect 199090 76650 199410 76850
rect 199480 76650 199520 76850
rect 199590 76650 199910 76850
rect 199980 76650 200020 76850
rect 200090 76650 200410 76850
rect 200480 76650 200520 76850
rect 200590 76650 200910 76850
rect 200980 76650 201020 76850
rect 201090 76650 201410 76850
rect 201480 76650 201520 76850
rect 201590 76650 201910 76850
rect 201980 76650 202020 76850
rect 202090 76650 202410 76850
rect 202480 76650 202520 76850
rect 202590 76650 202910 76850
rect 202980 76650 203020 76850
rect 203090 76650 203410 76850
rect 203480 76650 203520 76850
rect 203590 76650 203910 76850
rect 203980 76650 204020 76850
rect 204090 76650 204410 76850
rect 204480 76650 204520 76850
rect 204590 76650 204910 76850
rect 204980 76650 205020 76850
rect 205090 76650 205410 76850
rect 205480 76650 205520 76850
rect 205590 76650 205910 76850
rect 205980 76650 206020 76850
rect 206090 76650 206410 76850
rect 206480 76650 206520 76850
rect 206590 76650 206910 76850
rect 206980 76650 207020 76850
rect 207090 76650 207410 76850
rect 207480 76650 207520 76850
rect 207590 76650 207910 76850
rect 207980 76650 208000 76850
rect 196000 76640 208000 76650
rect 196140 76590 196360 76640
rect 196140 76520 196150 76590
rect 196350 76520 196360 76590
rect 196140 76480 196360 76520
rect 196140 76410 196150 76480
rect 196350 76410 196360 76480
rect 196140 76360 196360 76410
rect 196640 76590 196860 76640
rect 196640 76520 196650 76590
rect 196850 76520 196860 76590
rect 196640 76480 196860 76520
rect 196640 76410 196650 76480
rect 196850 76410 196860 76480
rect 196640 76360 196860 76410
rect 197140 76590 197360 76640
rect 197140 76520 197150 76590
rect 197350 76520 197360 76590
rect 197140 76480 197360 76520
rect 197140 76410 197150 76480
rect 197350 76410 197360 76480
rect 197140 76360 197360 76410
rect 197640 76590 197860 76640
rect 197640 76520 197650 76590
rect 197850 76520 197860 76590
rect 197640 76480 197860 76520
rect 197640 76410 197650 76480
rect 197850 76410 197860 76480
rect 197640 76360 197860 76410
rect 198140 76590 198360 76640
rect 198140 76520 198150 76590
rect 198350 76520 198360 76590
rect 198140 76480 198360 76520
rect 198140 76410 198150 76480
rect 198350 76410 198360 76480
rect 198140 76360 198360 76410
rect 198640 76590 198860 76640
rect 198640 76520 198650 76590
rect 198850 76520 198860 76590
rect 198640 76480 198860 76520
rect 198640 76410 198650 76480
rect 198850 76410 198860 76480
rect 198640 76360 198860 76410
rect 199140 76590 199360 76640
rect 199140 76520 199150 76590
rect 199350 76520 199360 76590
rect 199140 76480 199360 76520
rect 199140 76410 199150 76480
rect 199350 76410 199360 76480
rect 199140 76360 199360 76410
rect 199640 76590 199860 76640
rect 199640 76520 199650 76590
rect 199850 76520 199860 76590
rect 199640 76480 199860 76520
rect 199640 76410 199650 76480
rect 199850 76410 199860 76480
rect 199640 76360 199860 76410
rect 200140 76590 200360 76640
rect 200140 76520 200150 76590
rect 200350 76520 200360 76590
rect 200140 76480 200360 76520
rect 200140 76410 200150 76480
rect 200350 76410 200360 76480
rect 200140 76360 200360 76410
rect 200640 76590 200860 76640
rect 200640 76520 200650 76590
rect 200850 76520 200860 76590
rect 200640 76480 200860 76520
rect 200640 76410 200650 76480
rect 200850 76410 200860 76480
rect 200640 76360 200860 76410
rect 201140 76590 201360 76640
rect 201140 76520 201150 76590
rect 201350 76520 201360 76590
rect 201140 76480 201360 76520
rect 201140 76410 201150 76480
rect 201350 76410 201360 76480
rect 201140 76360 201360 76410
rect 201640 76590 201860 76640
rect 201640 76520 201650 76590
rect 201850 76520 201860 76590
rect 201640 76480 201860 76520
rect 201640 76410 201650 76480
rect 201850 76410 201860 76480
rect 201640 76360 201860 76410
rect 202140 76590 202360 76640
rect 202140 76520 202150 76590
rect 202350 76520 202360 76590
rect 202140 76480 202360 76520
rect 202140 76410 202150 76480
rect 202350 76410 202360 76480
rect 202140 76360 202360 76410
rect 202640 76590 202860 76640
rect 202640 76520 202650 76590
rect 202850 76520 202860 76590
rect 202640 76480 202860 76520
rect 202640 76410 202650 76480
rect 202850 76410 202860 76480
rect 202640 76360 202860 76410
rect 203140 76590 203360 76640
rect 203140 76520 203150 76590
rect 203350 76520 203360 76590
rect 203140 76480 203360 76520
rect 203140 76410 203150 76480
rect 203350 76410 203360 76480
rect 203140 76360 203360 76410
rect 203640 76590 203860 76640
rect 203640 76520 203650 76590
rect 203850 76520 203860 76590
rect 203640 76480 203860 76520
rect 203640 76410 203650 76480
rect 203850 76410 203860 76480
rect 203640 76360 203860 76410
rect 204140 76590 204360 76640
rect 204140 76520 204150 76590
rect 204350 76520 204360 76590
rect 204140 76480 204360 76520
rect 204140 76410 204150 76480
rect 204350 76410 204360 76480
rect 204140 76360 204360 76410
rect 204640 76590 204860 76640
rect 204640 76520 204650 76590
rect 204850 76520 204860 76590
rect 204640 76480 204860 76520
rect 204640 76410 204650 76480
rect 204850 76410 204860 76480
rect 204640 76360 204860 76410
rect 205140 76590 205360 76640
rect 205140 76520 205150 76590
rect 205350 76520 205360 76590
rect 205140 76480 205360 76520
rect 205140 76410 205150 76480
rect 205350 76410 205360 76480
rect 205140 76360 205360 76410
rect 205640 76590 205860 76640
rect 205640 76520 205650 76590
rect 205850 76520 205860 76590
rect 205640 76480 205860 76520
rect 205640 76410 205650 76480
rect 205850 76410 205860 76480
rect 205640 76360 205860 76410
rect 206140 76590 206360 76640
rect 206140 76520 206150 76590
rect 206350 76520 206360 76590
rect 206140 76480 206360 76520
rect 206140 76410 206150 76480
rect 206350 76410 206360 76480
rect 206140 76360 206360 76410
rect 206640 76590 206860 76640
rect 206640 76520 206650 76590
rect 206850 76520 206860 76590
rect 206640 76480 206860 76520
rect 206640 76410 206650 76480
rect 206850 76410 206860 76480
rect 206640 76360 206860 76410
rect 207140 76590 207360 76640
rect 207140 76520 207150 76590
rect 207350 76520 207360 76590
rect 207140 76480 207360 76520
rect 207140 76410 207150 76480
rect 207350 76410 207360 76480
rect 207140 76360 207360 76410
rect 207640 76590 207860 76640
rect 207640 76520 207650 76590
rect 207850 76520 207860 76590
rect 207640 76480 207860 76520
rect 207640 76410 207650 76480
rect 207850 76410 207860 76480
rect 207640 76360 207860 76410
rect 196000 76350 208000 76360
rect 196000 76150 196020 76350
rect 196090 76150 196410 76350
rect 196480 76150 196520 76350
rect 196590 76150 196910 76350
rect 196980 76150 197020 76350
rect 197090 76150 197410 76350
rect 197480 76150 197520 76350
rect 197590 76150 197910 76350
rect 197980 76150 198020 76350
rect 198090 76150 198410 76350
rect 198480 76150 198520 76350
rect 198590 76150 198910 76350
rect 198980 76150 199020 76350
rect 199090 76150 199410 76350
rect 199480 76150 199520 76350
rect 199590 76150 199910 76350
rect 199980 76150 200020 76350
rect 200090 76150 200410 76350
rect 200480 76150 200520 76350
rect 200590 76150 200910 76350
rect 200980 76150 201020 76350
rect 201090 76150 201410 76350
rect 201480 76150 201520 76350
rect 201590 76150 201910 76350
rect 201980 76150 202020 76350
rect 202090 76150 202410 76350
rect 202480 76150 202520 76350
rect 202590 76150 202910 76350
rect 202980 76150 203020 76350
rect 203090 76150 203410 76350
rect 203480 76150 203520 76350
rect 203590 76150 203910 76350
rect 203980 76150 204020 76350
rect 204090 76150 204410 76350
rect 204480 76150 204520 76350
rect 204590 76150 204910 76350
rect 204980 76150 205020 76350
rect 205090 76150 205410 76350
rect 205480 76150 205520 76350
rect 205590 76150 205910 76350
rect 205980 76150 206020 76350
rect 206090 76150 206410 76350
rect 206480 76150 206520 76350
rect 206590 76150 206910 76350
rect 206980 76150 207020 76350
rect 207090 76150 207410 76350
rect 207480 76150 207520 76350
rect 207590 76150 207910 76350
rect 207980 76150 208000 76350
rect 196000 76140 208000 76150
rect 196140 76090 196360 76140
rect 196140 76020 196150 76090
rect 196350 76020 196360 76090
rect 196140 75980 196360 76020
rect 196140 75910 196150 75980
rect 196350 75910 196360 75980
rect 196140 75860 196360 75910
rect 196640 76090 196860 76140
rect 196640 76020 196650 76090
rect 196850 76020 196860 76090
rect 196640 75980 196860 76020
rect 196640 75910 196650 75980
rect 196850 75910 196860 75980
rect 196640 75860 196860 75910
rect 197140 76090 197360 76140
rect 197140 76020 197150 76090
rect 197350 76020 197360 76090
rect 197140 75980 197360 76020
rect 197140 75910 197150 75980
rect 197350 75910 197360 75980
rect 197140 75860 197360 75910
rect 197640 76090 197860 76140
rect 197640 76020 197650 76090
rect 197850 76020 197860 76090
rect 197640 75980 197860 76020
rect 197640 75910 197650 75980
rect 197850 75910 197860 75980
rect 197640 75860 197860 75910
rect 198140 76090 198360 76140
rect 198140 76020 198150 76090
rect 198350 76020 198360 76090
rect 198140 75980 198360 76020
rect 198140 75910 198150 75980
rect 198350 75910 198360 75980
rect 198140 75860 198360 75910
rect 198640 76090 198860 76140
rect 198640 76020 198650 76090
rect 198850 76020 198860 76090
rect 198640 75980 198860 76020
rect 198640 75910 198650 75980
rect 198850 75910 198860 75980
rect 198640 75860 198860 75910
rect 199140 76090 199360 76140
rect 199140 76020 199150 76090
rect 199350 76020 199360 76090
rect 199140 75980 199360 76020
rect 199140 75910 199150 75980
rect 199350 75910 199360 75980
rect 199140 75860 199360 75910
rect 199640 76090 199860 76140
rect 199640 76020 199650 76090
rect 199850 76020 199860 76090
rect 199640 75980 199860 76020
rect 199640 75910 199650 75980
rect 199850 75910 199860 75980
rect 199640 75860 199860 75910
rect 200140 76090 200360 76140
rect 200140 76020 200150 76090
rect 200350 76020 200360 76090
rect 200140 75980 200360 76020
rect 200140 75910 200150 75980
rect 200350 75910 200360 75980
rect 200140 75860 200360 75910
rect 200640 76090 200860 76140
rect 200640 76020 200650 76090
rect 200850 76020 200860 76090
rect 200640 75980 200860 76020
rect 200640 75910 200650 75980
rect 200850 75910 200860 75980
rect 200640 75860 200860 75910
rect 201140 76090 201360 76140
rect 201140 76020 201150 76090
rect 201350 76020 201360 76090
rect 201140 75980 201360 76020
rect 201140 75910 201150 75980
rect 201350 75910 201360 75980
rect 201140 75860 201360 75910
rect 201640 76090 201860 76140
rect 201640 76020 201650 76090
rect 201850 76020 201860 76090
rect 201640 75980 201860 76020
rect 201640 75910 201650 75980
rect 201850 75910 201860 75980
rect 201640 75860 201860 75910
rect 202140 76090 202360 76140
rect 202140 76020 202150 76090
rect 202350 76020 202360 76090
rect 202140 75980 202360 76020
rect 202140 75910 202150 75980
rect 202350 75910 202360 75980
rect 202140 75860 202360 75910
rect 202640 76090 202860 76140
rect 202640 76020 202650 76090
rect 202850 76020 202860 76090
rect 202640 75980 202860 76020
rect 202640 75910 202650 75980
rect 202850 75910 202860 75980
rect 202640 75860 202860 75910
rect 203140 76090 203360 76140
rect 203140 76020 203150 76090
rect 203350 76020 203360 76090
rect 203140 75980 203360 76020
rect 203140 75910 203150 75980
rect 203350 75910 203360 75980
rect 203140 75860 203360 75910
rect 203640 76090 203860 76140
rect 203640 76020 203650 76090
rect 203850 76020 203860 76090
rect 203640 75980 203860 76020
rect 203640 75910 203650 75980
rect 203850 75910 203860 75980
rect 203640 75860 203860 75910
rect 204140 76090 204360 76140
rect 204140 76020 204150 76090
rect 204350 76020 204360 76090
rect 204140 75980 204360 76020
rect 204140 75910 204150 75980
rect 204350 75910 204360 75980
rect 204140 75860 204360 75910
rect 204640 76090 204860 76140
rect 204640 76020 204650 76090
rect 204850 76020 204860 76090
rect 204640 75980 204860 76020
rect 204640 75910 204650 75980
rect 204850 75910 204860 75980
rect 204640 75860 204860 75910
rect 205140 76090 205360 76140
rect 205140 76020 205150 76090
rect 205350 76020 205360 76090
rect 205140 75980 205360 76020
rect 205140 75910 205150 75980
rect 205350 75910 205360 75980
rect 205140 75860 205360 75910
rect 205640 76090 205860 76140
rect 205640 76020 205650 76090
rect 205850 76020 205860 76090
rect 205640 75980 205860 76020
rect 205640 75910 205650 75980
rect 205850 75910 205860 75980
rect 205640 75860 205860 75910
rect 206140 76090 206360 76140
rect 206140 76020 206150 76090
rect 206350 76020 206360 76090
rect 206140 75980 206360 76020
rect 206140 75910 206150 75980
rect 206350 75910 206360 75980
rect 206140 75860 206360 75910
rect 206640 76090 206860 76140
rect 206640 76020 206650 76090
rect 206850 76020 206860 76090
rect 206640 75980 206860 76020
rect 206640 75910 206650 75980
rect 206850 75910 206860 75980
rect 206640 75860 206860 75910
rect 207140 76090 207360 76140
rect 207140 76020 207150 76090
rect 207350 76020 207360 76090
rect 207140 75980 207360 76020
rect 207140 75910 207150 75980
rect 207350 75910 207360 75980
rect 207140 75860 207360 75910
rect 207640 76090 207860 76140
rect 207640 76020 207650 76090
rect 207850 76020 207860 76090
rect 207640 75980 207860 76020
rect 207640 75910 207650 75980
rect 207850 75910 207860 75980
rect 207640 75860 207860 75910
rect 196000 75850 208000 75860
rect 196000 75650 196020 75850
rect 196090 75650 196410 75850
rect 196480 75650 196520 75850
rect 196590 75650 196910 75850
rect 196980 75650 197020 75850
rect 197090 75650 197410 75850
rect 197480 75650 197520 75850
rect 197590 75650 197910 75850
rect 197980 75650 198020 75850
rect 198090 75650 198410 75850
rect 198480 75650 198520 75850
rect 198590 75650 198910 75850
rect 198980 75650 199020 75850
rect 199090 75650 199410 75850
rect 199480 75650 199520 75850
rect 199590 75650 199910 75850
rect 199980 75650 200020 75850
rect 200090 75650 200410 75850
rect 200480 75650 200520 75850
rect 200590 75650 200910 75850
rect 200980 75650 201020 75850
rect 201090 75650 201410 75850
rect 201480 75650 201520 75850
rect 201590 75650 201910 75850
rect 201980 75650 202020 75850
rect 202090 75650 202410 75850
rect 202480 75650 202520 75850
rect 202590 75650 202910 75850
rect 202980 75650 203020 75850
rect 203090 75650 203410 75850
rect 203480 75650 203520 75850
rect 203590 75650 203910 75850
rect 203980 75650 204020 75850
rect 204090 75650 204410 75850
rect 204480 75650 204520 75850
rect 204590 75650 204910 75850
rect 204980 75650 205020 75850
rect 205090 75650 205410 75850
rect 205480 75650 205520 75850
rect 205590 75650 205910 75850
rect 205980 75650 206020 75850
rect 206090 75650 206410 75850
rect 206480 75650 206520 75850
rect 206590 75650 206910 75850
rect 206980 75650 207020 75850
rect 207090 75650 207410 75850
rect 207480 75650 207520 75850
rect 207590 75650 207910 75850
rect 207980 75650 208000 75850
rect 196000 75640 208000 75650
rect 196140 75590 196360 75640
rect 196140 75520 196150 75590
rect 196350 75520 196360 75590
rect 196140 75480 196360 75520
rect 196140 75410 196150 75480
rect 196350 75410 196360 75480
rect 196140 75360 196360 75410
rect 196640 75590 196860 75640
rect 196640 75520 196650 75590
rect 196850 75520 196860 75590
rect 196640 75480 196860 75520
rect 196640 75410 196650 75480
rect 196850 75410 196860 75480
rect 196640 75360 196860 75410
rect 197140 75590 197360 75640
rect 197140 75520 197150 75590
rect 197350 75520 197360 75590
rect 197140 75480 197360 75520
rect 197140 75410 197150 75480
rect 197350 75410 197360 75480
rect 197140 75360 197360 75410
rect 197640 75590 197860 75640
rect 197640 75520 197650 75590
rect 197850 75520 197860 75590
rect 197640 75480 197860 75520
rect 197640 75410 197650 75480
rect 197850 75410 197860 75480
rect 197640 75360 197860 75410
rect 198140 75590 198360 75640
rect 198140 75520 198150 75590
rect 198350 75520 198360 75590
rect 198140 75480 198360 75520
rect 198140 75410 198150 75480
rect 198350 75410 198360 75480
rect 198140 75360 198360 75410
rect 198640 75590 198860 75640
rect 198640 75520 198650 75590
rect 198850 75520 198860 75590
rect 198640 75480 198860 75520
rect 198640 75410 198650 75480
rect 198850 75410 198860 75480
rect 198640 75360 198860 75410
rect 199140 75590 199360 75640
rect 199140 75520 199150 75590
rect 199350 75520 199360 75590
rect 199140 75480 199360 75520
rect 199140 75410 199150 75480
rect 199350 75410 199360 75480
rect 199140 75360 199360 75410
rect 199640 75590 199860 75640
rect 199640 75520 199650 75590
rect 199850 75520 199860 75590
rect 199640 75480 199860 75520
rect 199640 75410 199650 75480
rect 199850 75410 199860 75480
rect 199640 75360 199860 75410
rect 200140 75590 200360 75640
rect 200140 75520 200150 75590
rect 200350 75520 200360 75590
rect 200140 75480 200360 75520
rect 200140 75410 200150 75480
rect 200350 75410 200360 75480
rect 200140 75360 200360 75410
rect 200640 75590 200860 75640
rect 200640 75520 200650 75590
rect 200850 75520 200860 75590
rect 200640 75480 200860 75520
rect 200640 75410 200650 75480
rect 200850 75410 200860 75480
rect 200640 75360 200860 75410
rect 201140 75590 201360 75640
rect 201140 75520 201150 75590
rect 201350 75520 201360 75590
rect 201140 75480 201360 75520
rect 201140 75410 201150 75480
rect 201350 75410 201360 75480
rect 201140 75360 201360 75410
rect 201640 75590 201860 75640
rect 201640 75520 201650 75590
rect 201850 75520 201860 75590
rect 201640 75480 201860 75520
rect 201640 75410 201650 75480
rect 201850 75410 201860 75480
rect 201640 75360 201860 75410
rect 202140 75590 202360 75640
rect 202140 75520 202150 75590
rect 202350 75520 202360 75590
rect 202140 75480 202360 75520
rect 202140 75410 202150 75480
rect 202350 75410 202360 75480
rect 202140 75360 202360 75410
rect 202640 75590 202860 75640
rect 202640 75520 202650 75590
rect 202850 75520 202860 75590
rect 202640 75480 202860 75520
rect 202640 75410 202650 75480
rect 202850 75410 202860 75480
rect 202640 75360 202860 75410
rect 203140 75590 203360 75640
rect 203140 75520 203150 75590
rect 203350 75520 203360 75590
rect 203140 75480 203360 75520
rect 203140 75410 203150 75480
rect 203350 75410 203360 75480
rect 203140 75360 203360 75410
rect 203640 75590 203860 75640
rect 203640 75520 203650 75590
rect 203850 75520 203860 75590
rect 203640 75480 203860 75520
rect 203640 75410 203650 75480
rect 203850 75410 203860 75480
rect 203640 75360 203860 75410
rect 204140 75590 204360 75640
rect 204140 75520 204150 75590
rect 204350 75520 204360 75590
rect 204140 75480 204360 75520
rect 204140 75410 204150 75480
rect 204350 75410 204360 75480
rect 204140 75360 204360 75410
rect 204640 75590 204860 75640
rect 204640 75520 204650 75590
rect 204850 75520 204860 75590
rect 204640 75480 204860 75520
rect 204640 75410 204650 75480
rect 204850 75410 204860 75480
rect 204640 75360 204860 75410
rect 205140 75590 205360 75640
rect 205140 75520 205150 75590
rect 205350 75520 205360 75590
rect 205140 75480 205360 75520
rect 205140 75410 205150 75480
rect 205350 75410 205360 75480
rect 205140 75360 205360 75410
rect 205640 75590 205860 75640
rect 205640 75520 205650 75590
rect 205850 75520 205860 75590
rect 205640 75480 205860 75520
rect 205640 75410 205650 75480
rect 205850 75410 205860 75480
rect 205640 75360 205860 75410
rect 206140 75590 206360 75640
rect 206140 75520 206150 75590
rect 206350 75520 206360 75590
rect 206140 75480 206360 75520
rect 206140 75410 206150 75480
rect 206350 75410 206360 75480
rect 206140 75360 206360 75410
rect 206640 75590 206860 75640
rect 206640 75520 206650 75590
rect 206850 75520 206860 75590
rect 206640 75480 206860 75520
rect 206640 75410 206650 75480
rect 206850 75410 206860 75480
rect 206640 75360 206860 75410
rect 207140 75590 207360 75640
rect 207140 75520 207150 75590
rect 207350 75520 207360 75590
rect 207140 75480 207360 75520
rect 207140 75410 207150 75480
rect 207350 75410 207360 75480
rect 207140 75360 207360 75410
rect 207640 75590 207860 75640
rect 207640 75520 207650 75590
rect 207850 75520 207860 75590
rect 207640 75480 207860 75520
rect 207640 75410 207650 75480
rect 207850 75410 207860 75480
rect 207640 75360 207860 75410
rect 196000 75350 208000 75360
rect 196000 75150 196020 75350
rect 196090 75150 196410 75350
rect 196480 75150 196520 75350
rect 196590 75150 196910 75350
rect 196980 75150 197020 75350
rect 197090 75150 197410 75350
rect 197480 75150 197520 75350
rect 197590 75150 197910 75350
rect 197980 75150 198020 75350
rect 198090 75150 198410 75350
rect 198480 75150 198520 75350
rect 198590 75150 198910 75350
rect 198980 75150 199020 75350
rect 199090 75150 199410 75350
rect 199480 75150 199520 75350
rect 199590 75150 199910 75350
rect 199980 75150 200020 75350
rect 200090 75150 200410 75350
rect 200480 75150 200520 75350
rect 200590 75150 200910 75350
rect 200980 75150 201020 75350
rect 201090 75150 201410 75350
rect 201480 75150 201520 75350
rect 201590 75150 201910 75350
rect 201980 75150 202020 75350
rect 202090 75150 202410 75350
rect 202480 75150 202520 75350
rect 202590 75150 202910 75350
rect 202980 75150 203020 75350
rect 203090 75150 203410 75350
rect 203480 75150 203520 75350
rect 203590 75150 203910 75350
rect 203980 75150 204020 75350
rect 204090 75150 204410 75350
rect 204480 75150 204520 75350
rect 204590 75150 204910 75350
rect 204980 75150 205020 75350
rect 205090 75150 205410 75350
rect 205480 75150 205520 75350
rect 205590 75150 205910 75350
rect 205980 75150 206020 75350
rect 206090 75150 206410 75350
rect 206480 75150 206520 75350
rect 206590 75150 206910 75350
rect 206980 75150 207020 75350
rect 207090 75150 207410 75350
rect 207480 75150 207520 75350
rect 207590 75150 207910 75350
rect 207980 75150 208000 75350
rect 196000 75140 208000 75150
rect 196140 75090 196360 75140
rect 196140 75020 196150 75090
rect 196350 75020 196360 75090
rect 196140 74980 196360 75020
rect 196140 74910 196150 74980
rect 196350 74910 196360 74980
rect 196140 74860 196360 74910
rect 196640 75090 196860 75140
rect 196640 75020 196650 75090
rect 196850 75020 196860 75090
rect 196640 74980 196860 75020
rect 196640 74910 196650 74980
rect 196850 74910 196860 74980
rect 196640 74860 196860 74910
rect 197140 75090 197360 75140
rect 197140 75020 197150 75090
rect 197350 75020 197360 75090
rect 197140 74980 197360 75020
rect 197140 74910 197150 74980
rect 197350 74910 197360 74980
rect 197140 74860 197360 74910
rect 197640 75090 197860 75140
rect 197640 75020 197650 75090
rect 197850 75020 197860 75090
rect 197640 74980 197860 75020
rect 197640 74910 197650 74980
rect 197850 74910 197860 74980
rect 197640 74860 197860 74910
rect 198140 75090 198360 75140
rect 198140 75020 198150 75090
rect 198350 75020 198360 75090
rect 198140 74980 198360 75020
rect 198140 74910 198150 74980
rect 198350 74910 198360 74980
rect 198140 74860 198360 74910
rect 198640 75090 198860 75140
rect 198640 75020 198650 75090
rect 198850 75020 198860 75090
rect 198640 74980 198860 75020
rect 198640 74910 198650 74980
rect 198850 74910 198860 74980
rect 198640 74860 198860 74910
rect 199140 75090 199360 75140
rect 199140 75020 199150 75090
rect 199350 75020 199360 75090
rect 199140 74980 199360 75020
rect 199140 74910 199150 74980
rect 199350 74910 199360 74980
rect 199140 74860 199360 74910
rect 199640 75090 199860 75140
rect 199640 75020 199650 75090
rect 199850 75020 199860 75090
rect 199640 74980 199860 75020
rect 199640 74910 199650 74980
rect 199850 74910 199860 74980
rect 199640 74860 199860 74910
rect 200140 75090 200360 75140
rect 200140 75020 200150 75090
rect 200350 75020 200360 75090
rect 200140 74980 200360 75020
rect 200140 74910 200150 74980
rect 200350 74910 200360 74980
rect 200140 74860 200360 74910
rect 200640 75090 200860 75140
rect 200640 75020 200650 75090
rect 200850 75020 200860 75090
rect 200640 74980 200860 75020
rect 200640 74910 200650 74980
rect 200850 74910 200860 74980
rect 200640 74860 200860 74910
rect 201140 75090 201360 75140
rect 201140 75020 201150 75090
rect 201350 75020 201360 75090
rect 201140 74980 201360 75020
rect 201140 74910 201150 74980
rect 201350 74910 201360 74980
rect 201140 74860 201360 74910
rect 201640 75090 201860 75140
rect 201640 75020 201650 75090
rect 201850 75020 201860 75090
rect 201640 74980 201860 75020
rect 201640 74910 201650 74980
rect 201850 74910 201860 74980
rect 201640 74860 201860 74910
rect 202140 75090 202360 75140
rect 202140 75020 202150 75090
rect 202350 75020 202360 75090
rect 202140 74980 202360 75020
rect 202140 74910 202150 74980
rect 202350 74910 202360 74980
rect 202140 74860 202360 74910
rect 202640 75090 202860 75140
rect 202640 75020 202650 75090
rect 202850 75020 202860 75090
rect 202640 74980 202860 75020
rect 202640 74910 202650 74980
rect 202850 74910 202860 74980
rect 202640 74860 202860 74910
rect 203140 75090 203360 75140
rect 203140 75020 203150 75090
rect 203350 75020 203360 75090
rect 203140 74980 203360 75020
rect 203140 74910 203150 74980
rect 203350 74910 203360 74980
rect 203140 74860 203360 74910
rect 203640 75090 203860 75140
rect 203640 75020 203650 75090
rect 203850 75020 203860 75090
rect 203640 74980 203860 75020
rect 203640 74910 203650 74980
rect 203850 74910 203860 74980
rect 203640 74860 203860 74910
rect 204140 75090 204360 75140
rect 204140 75020 204150 75090
rect 204350 75020 204360 75090
rect 204140 74980 204360 75020
rect 204140 74910 204150 74980
rect 204350 74910 204360 74980
rect 204140 74860 204360 74910
rect 204640 75090 204860 75140
rect 204640 75020 204650 75090
rect 204850 75020 204860 75090
rect 204640 74980 204860 75020
rect 204640 74910 204650 74980
rect 204850 74910 204860 74980
rect 204640 74860 204860 74910
rect 205140 75090 205360 75140
rect 205140 75020 205150 75090
rect 205350 75020 205360 75090
rect 205140 74980 205360 75020
rect 205140 74910 205150 74980
rect 205350 74910 205360 74980
rect 205140 74860 205360 74910
rect 205640 75090 205860 75140
rect 205640 75020 205650 75090
rect 205850 75020 205860 75090
rect 205640 74980 205860 75020
rect 205640 74910 205650 74980
rect 205850 74910 205860 74980
rect 205640 74860 205860 74910
rect 206140 75090 206360 75140
rect 206140 75020 206150 75090
rect 206350 75020 206360 75090
rect 206140 74980 206360 75020
rect 206140 74910 206150 74980
rect 206350 74910 206360 74980
rect 206140 74860 206360 74910
rect 206640 75090 206860 75140
rect 206640 75020 206650 75090
rect 206850 75020 206860 75090
rect 206640 74980 206860 75020
rect 206640 74910 206650 74980
rect 206850 74910 206860 74980
rect 206640 74860 206860 74910
rect 207140 75090 207360 75140
rect 207140 75020 207150 75090
rect 207350 75020 207360 75090
rect 207140 74980 207360 75020
rect 207140 74910 207150 74980
rect 207350 74910 207360 74980
rect 207140 74860 207360 74910
rect 207640 75090 207860 75140
rect 207640 75020 207650 75090
rect 207850 75020 207860 75090
rect 207640 74980 207860 75020
rect 207640 74910 207650 74980
rect 207850 74910 207860 74980
rect 207640 74860 207860 74910
rect 196000 74850 208000 74860
rect 196000 74650 196020 74850
rect 196090 74650 196410 74850
rect 196480 74650 196520 74850
rect 196590 74650 196910 74850
rect 196980 74650 197020 74850
rect 197090 74650 197410 74850
rect 197480 74650 197520 74850
rect 197590 74650 197910 74850
rect 197980 74650 198020 74850
rect 198090 74650 198410 74850
rect 198480 74650 198520 74850
rect 198590 74650 198910 74850
rect 198980 74650 199020 74850
rect 199090 74650 199410 74850
rect 199480 74650 199520 74850
rect 199590 74650 199910 74850
rect 199980 74650 200020 74850
rect 200090 74650 200410 74850
rect 200480 74650 200520 74850
rect 200590 74650 200910 74850
rect 200980 74650 201020 74850
rect 201090 74650 201410 74850
rect 201480 74650 201520 74850
rect 201590 74650 201910 74850
rect 201980 74650 202020 74850
rect 202090 74650 202410 74850
rect 202480 74650 202520 74850
rect 202590 74650 202910 74850
rect 202980 74650 203020 74850
rect 203090 74650 203410 74850
rect 203480 74650 203520 74850
rect 203590 74650 203910 74850
rect 203980 74650 204020 74850
rect 204090 74650 204410 74850
rect 204480 74650 204520 74850
rect 204590 74650 204910 74850
rect 204980 74650 205020 74850
rect 205090 74650 205410 74850
rect 205480 74650 205520 74850
rect 205590 74650 205910 74850
rect 205980 74650 206020 74850
rect 206090 74650 206410 74850
rect 206480 74650 206520 74850
rect 206590 74650 206910 74850
rect 206980 74650 207020 74850
rect 207090 74650 207410 74850
rect 207480 74650 207520 74850
rect 207590 74650 207910 74850
rect 207980 74650 208000 74850
rect 196000 74640 208000 74650
rect 196140 74590 196360 74640
rect 196140 74520 196150 74590
rect 196350 74520 196360 74590
rect 196140 74480 196360 74520
rect 196140 74410 196150 74480
rect 196350 74410 196360 74480
rect 196140 74360 196360 74410
rect 196640 74590 196860 74640
rect 196640 74520 196650 74590
rect 196850 74520 196860 74590
rect 196640 74480 196860 74520
rect 196640 74410 196650 74480
rect 196850 74410 196860 74480
rect 196640 74360 196860 74410
rect 197140 74590 197360 74640
rect 197140 74520 197150 74590
rect 197350 74520 197360 74590
rect 197140 74480 197360 74520
rect 197140 74410 197150 74480
rect 197350 74410 197360 74480
rect 197140 74360 197360 74410
rect 197640 74590 197860 74640
rect 197640 74520 197650 74590
rect 197850 74520 197860 74590
rect 197640 74480 197860 74520
rect 197640 74410 197650 74480
rect 197850 74410 197860 74480
rect 197640 74360 197860 74410
rect 198140 74590 198360 74640
rect 198140 74520 198150 74590
rect 198350 74520 198360 74590
rect 198140 74480 198360 74520
rect 198140 74410 198150 74480
rect 198350 74410 198360 74480
rect 198140 74360 198360 74410
rect 198640 74590 198860 74640
rect 198640 74520 198650 74590
rect 198850 74520 198860 74590
rect 198640 74480 198860 74520
rect 198640 74410 198650 74480
rect 198850 74410 198860 74480
rect 198640 74360 198860 74410
rect 199140 74590 199360 74640
rect 199140 74520 199150 74590
rect 199350 74520 199360 74590
rect 199140 74480 199360 74520
rect 199140 74410 199150 74480
rect 199350 74410 199360 74480
rect 199140 74360 199360 74410
rect 199640 74590 199860 74640
rect 199640 74520 199650 74590
rect 199850 74520 199860 74590
rect 199640 74480 199860 74520
rect 199640 74410 199650 74480
rect 199850 74410 199860 74480
rect 199640 74360 199860 74410
rect 200140 74590 200360 74640
rect 200140 74520 200150 74590
rect 200350 74520 200360 74590
rect 200140 74480 200360 74520
rect 200140 74410 200150 74480
rect 200350 74410 200360 74480
rect 200140 74360 200360 74410
rect 200640 74590 200860 74640
rect 200640 74520 200650 74590
rect 200850 74520 200860 74590
rect 200640 74480 200860 74520
rect 200640 74410 200650 74480
rect 200850 74410 200860 74480
rect 200640 74360 200860 74410
rect 201140 74590 201360 74640
rect 201140 74520 201150 74590
rect 201350 74520 201360 74590
rect 201140 74480 201360 74520
rect 201140 74410 201150 74480
rect 201350 74410 201360 74480
rect 201140 74360 201360 74410
rect 201640 74590 201860 74640
rect 201640 74520 201650 74590
rect 201850 74520 201860 74590
rect 201640 74480 201860 74520
rect 201640 74410 201650 74480
rect 201850 74410 201860 74480
rect 201640 74360 201860 74410
rect 202140 74590 202360 74640
rect 202140 74520 202150 74590
rect 202350 74520 202360 74590
rect 202140 74480 202360 74520
rect 202140 74410 202150 74480
rect 202350 74410 202360 74480
rect 202140 74360 202360 74410
rect 202640 74590 202860 74640
rect 202640 74520 202650 74590
rect 202850 74520 202860 74590
rect 202640 74480 202860 74520
rect 202640 74410 202650 74480
rect 202850 74410 202860 74480
rect 202640 74360 202860 74410
rect 203140 74590 203360 74640
rect 203140 74520 203150 74590
rect 203350 74520 203360 74590
rect 203140 74480 203360 74520
rect 203140 74410 203150 74480
rect 203350 74410 203360 74480
rect 203140 74360 203360 74410
rect 203640 74590 203860 74640
rect 203640 74520 203650 74590
rect 203850 74520 203860 74590
rect 203640 74480 203860 74520
rect 203640 74410 203650 74480
rect 203850 74410 203860 74480
rect 203640 74360 203860 74410
rect 204140 74590 204360 74640
rect 204140 74520 204150 74590
rect 204350 74520 204360 74590
rect 204140 74480 204360 74520
rect 204140 74410 204150 74480
rect 204350 74410 204360 74480
rect 204140 74360 204360 74410
rect 204640 74590 204860 74640
rect 204640 74520 204650 74590
rect 204850 74520 204860 74590
rect 204640 74480 204860 74520
rect 204640 74410 204650 74480
rect 204850 74410 204860 74480
rect 204640 74360 204860 74410
rect 205140 74590 205360 74640
rect 205140 74520 205150 74590
rect 205350 74520 205360 74590
rect 205140 74480 205360 74520
rect 205140 74410 205150 74480
rect 205350 74410 205360 74480
rect 205140 74360 205360 74410
rect 205640 74590 205860 74640
rect 205640 74520 205650 74590
rect 205850 74520 205860 74590
rect 205640 74480 205860 74520
rect 205640 74410 205650 74480
rect 205850 74410 205860 74480
rect 205640 74360 205860 74410
rect 206140 74590 206360 74640
rect 206140 74520 206150 74590
rect 206350 74520 206360 74590
rect 206140 74480 206360 74520
rect 206140 74410 206150 74480
rect 206350 74410 206360 74480
rect 206140 74360 206360 74410
rect 206640 74590 206860 74640
rect 206640 74520 206650 74590
rect 206850 74520 206860 74590
rect 206640 74480 206860 74520
rect 206640 74410 206650 74480
rect 206850 74410 206860 74480
rect 206640 74360 206860 74410
rect 207140 74590 207360 74640
rect 207140 74520 207150 74590
rect 207350 74520 207360 74590
rect 207140 74480 207360 74520
rect 207140 74410 207150 74480
rect 207350 74410 207360 74480
rect 207140 74360 207360 74410
rect 207640 74590 207860 74640
rect 207640 74520 207650 74590
rect 207850 74520 207860 74590
rect 207640 74480 207860 74520
rect 207640 74410 207650 74480
rect 207850 74410 207860 74480
rect 207640 74360 207860 74410
rect 196000 74350 208000 74360
rect 196000 74150 196020 74350
rect 196090 74150 196410 74350
rect 196480 74150 196520 74350
rect 196590 74150 196910 74350
rect 196980 74150 197020 74350
rect 197090 74150 197410 74350
rect 197480 74150 197520 74350
rect 197590 74150 197910 74350
rect 197980 74150 198020 74350
rect 198090 74150 198410 74350
rect 198480 74150 198520 74350
rect 198590 74150 198910 74350
rect 198980 74150 199020 74350
rect 199090 74150 199410 74350
rect 199480 74150 199520 74350
rect 199590 74150 199910 74350
rect 199980 74150 200020 74350
rect 200090 74150 200410 74350
rect 200480 74150 200520 74350
rect 200590 74150 200910 74350
rect 200980 74150 201020 74350
rect 201090 74150 201410 74350
rect 201480 74150 201520 74350
rect 201590 74150 201910 74350
rect 201980 74150 202020 74350
rect 202090 74150 202410 74350
rect 202480 74150 202520 74350
rect 202590 74150 202910 74350
rect 202980 74150 203020 74350
rect 203090 74150 203410 74350
rect 203480 74150 203520 74350
rect 203590 74150 203910 74350
rect 203980 74150 204020 74350
rect 204090 74150 204410 74350
rect 204480 74150 204520 74350
rect 204590 74150 204910 74350
rect 204980 74150 205020 74350
rect 205090 74150 205410 74350
rect 205480 74150 205520 74350
rect 205590 74150 205910 74350
rect 205980 74150 206020 74350
rect 206090 74150 206410 74350
rect 206480 74150 206520 74350
rect 206590 74150 206910 74350
rect 206980 74150 207020 74350
rect 207090 74150 207410 74350
rect 207480 74150 207520 74350
rect 207590 74150 207910 74350
rect 207980 74150 208000 74350
rect 196000 74140 208000 74150
rect 196140 74090 196360 74140
rect 196140 74020 196150 74090
rect 196350 74020 196360 74090
rect 196140 73980 196360 74020
rect 196140 73910 196150 73980
rect 196350 73910 196360 73980
rect 196140 73860 196360 73910
rect 196640 74090 196860 74140
rect 196640 74020 196650 74090
rect 196850 74020 196860 74090
rect 196640 73980 196860 74020
rect 196640 73910 196650 73980
rect 196850 73910 196860 73980
rect 196640 73860 196860 73910
rect 197140 74090 197360 74140
rect 197140 74020 197150 74090
rect 197350 74020 197360 74090
rect 197140 73980 197360 74020
rect 197140 73910 197150 73980
rect 197350 73910 197360 73980
rect 197140 73860 197360 73910
rect 197640 74090 197860 74140
rect 197640 74020 197650 74090
rect 197850 74020 197860 74090
rect 197640 73980 197860 74020
rect 197640 73910 197650 73980
rect 197850 73910 197860 73980
rect 197640 73860 197860 73910
rect 198140 74090 198360 74140
rect 198140 74020 198150 74090
rect 198350 74020 198360 74090
rect 198140 73980 198360 74020
rect 198140 73910 198150 73980
rect 198350 73910 198360 73980
rect 198140 73860 198360 73910
rect 198640 74090 198860 74140
rect 198640 74020 198650 74090
rect 198850 74020 198860 74090
rect 198640 73980 198860 74020
rect 198640 73910 198650 73980
rect 198850 73910 198860 73980
rect 198640 73860 198860 73910
rect 199140 74090 199360 74140
rect 199140 74020 199150 74090
rect 199350 74020 199360 74090
rect 199140 73980 199360 74020
rect 199140 73910 199150 73980
rect 199350 73910 199360 73980
rect 199140 73860 199360 73910
rect 199640 74090 199860 74140
rect 199640 74020 199650 74090
rect 199850 74020 199860 74090
rect 199640 73980 199860 74020
rect 199640 73910 199650 73980
rect 199850 73910 199860 73980
rect 199640 73860 199860 73910
rect 200140 74090 200360 74140
rect 200140 74020 200150 74090
rect 200350 74020 200360 74090
rect 200140 73980 200360 74020
rect 200140 73910 200150 73980
rect 200350 73910 200360 73980
rect 200140 73860 200360 73910
rect 200640 74090 200860 74140
rect 200640 74020 200650 74090
rect 200850 74020 200860 74090
rect 200640 73980 200860 74020
rect 200640 73910 200650 73980
rect 200850 73910 200860 73980
rect 200640 73860 200860 73910
rect 201140 74090 201360 74140
rect 201140 74020 201150 74090
rect 201350 74020 201360 74090
rect 201140 73980 201360 74020
rect 201140 73910 201150 73980
rect 201350 73910 201360 73980
rect 201140 73860 201360 73910
rect 201640 74090 201860 74140
rect 201640 74020 201650 74090
rect 201850 74020 201860 74090
rect 201640 73980 201860 74020
rect 201640 73910 201650 73980
rect 201850 73910 201860 73980
rect 201640 73860 201860 73910
rect 202140 74090 202360 74140
rect 202140 74020 202150 74090
rect 202350 74020 202360 74090
rect 202140 73980 202360 74020
rect 202140 73910 202150 73980
rect 202350 73910 202360 73980
rect 202140 73860 202360 73910
rect 202640 74090 202860 74140
rect 202640 74020 202650 74090
rect 202850 74020 202860 74090
rect 202640 73980 202860 74020
rect 202640 73910 202650 73980
rect 202850 73910 202860 73980
rect 202640 73860 202860 73910
rect 203140 74090 203360 74140
rect 203140 74020 203150 74090
rect 203350 74020 203360 74090
rect 203140 73980 203360 74020
rect 203140 73910 203150 73980
rect 203350 73910 203360 73980
rect 203140 73860 203360 73910
rect 203640 74090 203860 74140
rect 203640 74020 203650 74090
rect 203850 74020 203860 74090
rect 203640 73980 203860 74020
rect 203640 73910 203650 73980
rect 203850 73910 203860 73980
rect 203640 73860 203860 73910
rect 204140 74090 204360 74140
rect 204140 74020 204150 74090
rect 204350 74020 204360 74090
rect 204140 73980 204360 74020
rect 204140 73910 204150 73980
rect 204350 73910 204360 73980
rect 204140 73860 204360 73910
rect 204640 74090 204860 74140
rect 204640 74020 204650 74090
rect 204850 74020 204860 74090
rect 204640 73980 204860 74020
rect 204640 73910 204650 73980
rect 204850 73910 204860 73980
rect 204640 73860 204860 73910
rect 205140 74090 205360 74140
rect 205140 74020 205150 74090
rect 205350 74020 205360 74090
rect 205140 73980 205360 74020
rect 205140 73910 205150 73980
rect 205350 73910 205360 73980
rect 205140 73860 205360 73910
rect 205640 74090 205860 74140
rect 205640 74020 205650 74090
rect 205850 74020 205860 74090
rect 205640 73980 205860 74020
rect 205640 73910 205650 73980
rect 205850 73910 205860 73980
rect 205640 73860 205860 73910
rect 206140 74090 206360 74140
rect 206140 74020 206150 74090
rect 206350 74020 206360 74090
rect 206140 73980 206360 74020
rect 206140 73910 206150 73980
rect 206350 73910 206360 73980
rect 206140 73860 206360 73910
rect 206640 74090 206860 74140
rect 206640 74020 206650 74090
rect 206850 74020 206860 74090
rect 206640 73980 206860 74020
rect 206640 73910 206650 73980
rect 206850 73910 206860 73980
rect 206640 73860 206860 73910
rect 207140 74090 207360 74140
rect 207140 74020 207150 74090
rect 207350 74020 207360 74090
rect 207140 73980 207360 74020
rect 207140 73910 207150 73980
rect 207350 73910 207360 73980
rect 207140 73860 207360 73910
rect 207640 74090 207860 74140
rect 207640 74020 207650 74090
rect 207850 74020 207860 74090
rect 207640 73980 207860 74020
rect 207640 73910 207650 73980
rect 207850 73910 207860 73980
rect 207640 73860 207860 73910
rect 196000 73850 208000 73860
rect 196000 73650 196020 73850
rect 196090 73650 196410 73850
rect 196480 73650 196520 73850
rect 196590 73650 196910 73850
rect 196980 73650 197020 73850
rect 197090 73650 197410 73850
rect 197480 73650 197520 73850
rect 197590 73650 197910 73850
rect 197980 73650 198020 73850
rect 198090 73650 198410 73850
rect 198480 73650 198520 73850
rect 198590 73650 198910 73850
rect 198980 73650 199020 73850
rect 199090 73650 199410 73850
rect 199480 73650 199520 73850
rect 199590 73650 199910 73850
rect 199980 73650 200020 73850
rect 200090 73650 200410 73850
rect 200480 73650 200520 73850
rect 200590 73650 200910 73850
rect 200980 73650 201020 73850
rect 201090 73650 201410 73850
rect 201480 73650 201520 73850
rect 201590 73650 201910 73850
rect 201980 73650 202020 73850
rect 202090 73650 202410 73850
rect 202480 73650 202520 73850
rect 202590 73650 202910 73850
rect 202980 73650 203020 73850
rect 203090 73650 203410 73850
rect 203480 73650 203520 73850
rect 203590 73650 203910 73850
rect 203980 73650 204020 73850
rect 204090 73650 204410 73850
rect 204480 73650 204520 73850
rect 204590 73650 204910 73850
rect 204980 73650 205020 73850
rect 205090 73650 205410 73850
rect 205480 73650 205520 73850
rect 205590 73650 205910 73850
rect 205980 73650 206020 73850
rect 206090 73650 206410 73850
rect 206480 73650 206520 73850
rect 206590 73650 206910 73850
rect 206980 73650 207020 73850
rect 207090 73650 207410 73850
rect 207480 73650 207520 73850
rect 207590 73650 207910 73850
rect 207980 73650 208000 73850
rect 196000 73640 208000 73650
rect 196140 73590 196360 73640
rect 196140 73520 196150 73590
rect 196350 73520 196360 73590
rect 196140 73480 196360 73520
rect 196140 73410 196150 73480
rect 196350 73410 196360 73480
rect 196140 73360 196360 73410
rect 196640 73590 196860 73640
rect 196640 73520 196650 73590
rect 196850 73520 196860 73590
rect 196640 73480 196860 73520
rect 196640 73410 196650 73480
rect 196850 73410 196860 73480
rect 196640 73360 196860 73410
rect 197140 73590 197360 73640
rect 197140 73520 197150 73590
rect 197350 73520 197360 73590
rect 197140 73480 197360 73520
rect 197140 73410 197150 73480
rect 197350 73410 197360 73480
rect 197140 73360 197360 73410
rect 197640 73590 197860 73640
rect 197640 73520 197650 73590
rect 197850 73520 197860 73590
rect 197640 73480 197860 73520
rect 197640 73410 197650 73480
rect 197850 73410 197860 73480
rect 197640 73360 197860 73410
rect 198140 73590 198360 73640
rect 198140 73520 198150 73590
rect 198350 73520 198360 73590
rect 198140 73480 198360 73520
rect 198140 73410 198150 73480
rect 198350 73410 198360 73480
rect 198140 73360 198360 73410
rect 198640 73590 198860 73640
rect 198640 73520 198650 73590
rect 198850 73520 198860 73590
rect 198640 73480 198860 73520
rect 198640 73410 198650 73480
rect 198850 73410 198860 73480
rect 198640 73360 198860 73410
rect 199140 73590 199360 73640
rect 199140 73520 199150 73590
rect 199350 73520 199360 73590
rect 199140 73480 199360 73520
rect 199140 73410 199150 73480
rect 199350 73410 199360 73480
rect 199140 73360 199360 73410
rect 199640 73590 199860 73640
rect 199640 73520 199650 73590
rect 199850 73520 199860 73590
rect 199640 73480 199860 73520
rect 199640 73410 199650 73480
rect 199850 73410 199860 73480
rect 199640 73360 199860 73410
rect 200140 73590 200360 73640
rect 200140 73520 200150 73590
rect 200350 73520 200360 73590
rect 200140 73480 200360 73520
rect 200140 73410 200150 73480
rect 200350 73410 200360 73480
rect 200140 73360 200360 73410
rect 200640 73590 200860 73640
rect 200640 73520 200650 73590
rect 200850 73520 200860 73590
rect 200640 73480 200860 73520
rect 200640 73410 200650 73480
rect 200850 73410 200860 73480
rect 200640 73360 200860 73410
rect 201140 73590 201360 73640
rect 201140 73520 201150 73590
rect 201350 73520 201360 73590
rect 201140 73480 201360 73520
rect 201140 73410 201150 73480
rect 201350 73410 201360 73480
rect 201140 73360 201360 73410
rect 201640 73590 201860 73640
rect 201640 73520 201650 73590
rect 201850 73520 201860 73590
rect 201640 73480 201860 73520
rect 201640 73410 201650 73480
rect 201850 73410 201860 73480
rect 201640 73360 201860 73410
rect 202140 73590 202360 73640
rect 202140 73520 202150 73590
rect 202350 73520 202360 73590
rect 202140 73480 202360 73520
rect 202140 73410 202150 73480
rect 202350 73410 202360 73480
rect 202140 73360 202360 73410
rect 202640 73590 202860 73640
rect 202640 73520 202650 73590
rect 202850 73520 202860 73590
rect 202640 73480 202860 73520
rect 202640 73410 202650 73480
rect 202850 73410 202860 73480
rect 202640 73360 202860 73410
rect 203140 73590 203360 73640
rect 203140 73520 203150 73590
rect 203350 73520 203360 73590
rect 203140 73480 203360 73520
rect 203140 73410 203150 73480
rect 203350 73410 203360 73480
rect 203140 73360 203360 73410
rect 203640 73590 203860 73640
rect 203640 73520 203650 73590
rect 203850 73520 203860 73590
rect 203640 73480 203860 73520
rect 203640 73410 203650 73480
rect 203850 73410 203860 73480
rect 203640 73360 203860 73410
rect 204140 73590 204360 73640
rect 204140 73520 204150 73590
rect 204350 73520 204360 73590
rect 204140 73480 204360 73520
rect 204140 73410 204150 73480
rect 204350 73410 204360 73480
rect 204140 73360 204360 73410
rect 204640 73590 204860 73640
rect 204640 73520 204650 73590
rect 204850 73520 204860 73590
rect 204640 73480 204860 73520
rect 204640 73410 204650 73480
rect 204850 73410 204860 73480
rect 204640 73360 204860 73410
rect 205140 73590 205360 73640
rect 205140 73520 205150 73590
rect 205350 73520 205360 73590
rect 205140 73480 205360 73520
rect 205140 73410 205150 73480
rect 205350 73410 205360 73480
rect 205140 73360 205360 73410
rect 205640 73590 205860 73640
rect 205640 73520 205650 73590
rect 205850 73520 205860 73590
rect 205640 73480 205860 73520
rect 205640 73410 205650 73480
rect 205850 73410 205860 73480
rect 205640 73360 205860 73410
rect 206140 73590 206360 73640
rect 206140 73520 206150 73590
rect 206350 73520 206360 73590
rect 206140 73480 206360 73520
rect 206140 73410 206150 73480
rect 206350 73410 206360 73480
rect 206140 73360 206360 73410
rect 206640 73590 206860 73640
rect 206640 73520 206650 73590
rect 206850 73520 206860 73590
rect 206640 73480 206860 73520
rect 206640 73410 206650 73480
rect 206850 73410 206860 73480
rect 206640 73360 206860 73410
rect 207140 73590 207360 73640
rect 207140 73520 207150 73590
rect 207350 73520 207360 73590
rect 207140 73480 207360 73520
rect 207140 73410 207150 73480
rect 207350 73410 207360 73480
rect 207140 73360 207360 73410
rect 207640 73590 207860 73640
rect 207640 73520 207650 73590
rect 207850 73520 207860 73590
rect 207640 73480 207860 73520
rect 207640 73410 207650 73480
rect 207850 73410 207860 73480
rect 207640 73360 207860 73410
rect 196000 73350 208000 73360
rect 196000 73150 196020 73350
rect 196090 73150 196410 73350
rect 196480 73150 196520 73350
rect 196590 73150 196910 73350
rect 196980 73150 197020 73350
rect 197090 73150 197410 73350
rect 197480 73150 197520 73350
rect 197590 73150 197910 73350
rect 197980 73150 198020 73350
rect 198090 73150 198410 73350
rect 198480 73150 198520 73350
rect 198590 73150 198910 73350
rect 198980 73150 199020 73350
rect 199090 73150 199410 73350
rect 199480 73150 199520 73350
rect 199590 73150 199910 73350
rect 199980 73150 200020 73350
rect 200090 73150 200410 73350
rect 200480 73150 200520 73350
rect 200590 73150 200910 73350
rect 200980 73150 201020 73350
rect 201090 73150 201410 73350
rect 201480 73150 201520 73350
rect 201590 73150 201910 73350
rect 201980 73150 202020 73350
rect 202090 73150 202410 73350
rect 202480 73150 202520 73350
rect 202590 73150 202910 73350
rect 202980 73150 203020 73350
rect 203090 73150 203410 73350
rect 203480 73150 203520 73350
rect 203590 73150 203910 73350
rect 203980 73150 204020 73350
rect 204090 73150 204410 73350
rect 204480 73150 204520 73350
rect 204590 73150 204910 73350
rect 204980 73150 205020 73350
rect 205090 73150 205410 73350
rect 205480 73150 205520 73350
rect 205590 73150 205910 73350
rect 205980 73150 206020 73350
rect 206090 73150 206410 73350
rect 206480 73150 206520 73350
rect 206590 73150 206910 73350
rect 206980 73150 207020 73350
rect 207090 73150 207410 73350
rect 207480 73150 207520 73350
rect 207590 73150 207910 73350
rect 207980 73150 208000 73350
rect 196000 73140 208000 73150
rect 196140 73090 196360 73140
rect 196140 73020 196150 73090
rect 196350 73020 196360 73090
rect 196140 72980 196360 73020
rect 196140 72910 196150 72980
rect 196350 72910 196360 72980
rect 196140 72860 196360 72910
rect 196640 73090 196860 73140
rect 196640 73020 196650 73090
rect 196850 73020 196860 73090
rect 196640 72980 196860 73020
rect 196640 72910 196650 72980
rect 196850 72910 196860 72980
rect 196640 72860 196860 72910
rect 197140 73090 197360 73140
rect 197140 73020 197150 73090
rect 197350 73020 197360 73090
rect 197140 72980 197360 73020
rect 197140 72910 197150 72980
rect 197350 72910 197360 72980
rect 197140 72860 197360 72910
rect 197640 73090 197860 73140
rect 197640 73020 197650 73090
rect 197850 73020 197860 73090
rect 197640 72980 197860 73020
rect 197640 72910 197650 72980
rect 197850 72910 197860 72980
rect 197640 72860 197860 72910
rect 198140 73090 198360 73140
rect 198140 73020 198150 73090
rect 198350 73020 198360 73090
rect 198140 72980 198360 73020
rect 198140 72910 198150 72980
rect 198350 72910 198360 72980
rect 198140 72860 198360 72910
rect 198640 73090 198860 73140
rect 198640 73020 198650 73090
rect 198850 73020 198860 73090
rect 198640 72980 198860 73020
rect 198640 72910 198650 72980
rect 198850 72910 198860 72980
rect 198640 72860 198860 72910
rect 199140 73090 199360 73140
rect 199140 73020 199150 73090
rect 199350 73020 199360 73090
rect 199140 72980 199360 73020
rect 199140 72910 199150 72980
rect 199350 72910 199360 72980
rect 199140 72860 199360 72910
rect 199640 73090 199860 73140
rect 199640 73020 199650 73090
rect 199850 73020 199860 73090
rect 199640 72980 199860 73020
rect 199640 72910 199650 72980
rect 199850 72910 199860 72980
rect 199640 72860 199860 72910
rect 200140 73090 200360 73140
rect 200140 73020 200150 73090
rect 200350 73020 200360 73090
rect 200140 72980 200360 73020
rect 200140 72910 200150 72980
rect 200350 72910 200360 72980
rect 200140 72860 200360 72910
rect 200640 73090 200860 73140
rect 200640 73020 200650 73090
rect 200850 73020 200860 73090
rect 200640 72980 200860 73020
rect 200640 72910 200650 72980
rect 200850 72910 200860 72980
rect 200640 72860 200860 72910
rect 201140 73090 201360 73140
rect 201140 73020 201150 73090
rect 201350 73020 201360 73090
rect 201140 72980 201360 73020
rect 201140 72910 201150 72980
rect 201350 72910 201360 72980
rect 201140 72860 201360 72910
rect 201640 73090 201860 73140
rect 201640 73020 201650 73090
rect 201850 73020 201860 73090
rect 201640 72980 201860 73020
rect 201640 72910 201650 72980
rect 201850 72910 201860 72980
rect 201640 72860 201860 72910
rect 202140 73090 202360 73140
rect 202140 73020 202150 73090
rect 202350 73020 202360 73090
rect 202140 72980 202360 73020
rect 202140 72910 202150 72980
rect 202350 72910 202360 72980
rect 202140 72860 202360 72910
rect 202640 73090 202860 73140
rect 202640 73020 202650 73090
rect 202850 73020 202860 73090
rect 202640 72980 202860 73020
rect 202640 72910 202650 72980
rect 202850 72910 202860 72980
rect 202640 72860 202860 72910
rect 203140 73090 203360 73140
rect 203140 73020 203150 73090
rect 203350 73020 203360 73090
rect 203140 72980 203360 73020
rect 203140 72910 203150 72980
rect 203350 72910 203360 72980
rect 203140 72860 203360 72910
rect 203640 73090 203860 73140
rect 203640 73020 203650 73090
rect 203850 73020 203860 73090
rect 203640 72980 203860 73020
rect 203640 72910 203650 72980
rect 203850 72910 203860 72980
rect 203640 72860 203860 72910
rect 204140 73090 204360 73140
rect 204140 73020 204150 73090
rect 204350 73020 204360 73090
rect 204140 72980 204360 73020
rect 204140 72910 204150 72980
rect 204350 72910 204360 72980
rect 204140 72860 204360 72910
rect 204640 73090 204860 73140
rect 204640 73020 204650 73090
rect 204850 73020 204860 73090
rect 204640 72980 204860 73020
rect 204640 72910 204650 72980
rect 204850 72910 204860 72980
rect 204640 72860 204860 72910
rect 205140 73090 205360 73140
rect 205140 73020 205150 73090
rect 205350 73020 205360 73090
rect 205140 72980 205360 73020
rect 205140 72910 205150 72980
rect 205350 72910 205360 72980
rect 205140 72860 205360 72910
rect 205640 73090 205860 73140
rect 205640 73020 205650 73090
rect 205850 73020 205860 73090
rect 205640 72980 205860 73020
rect 205640 72910 205650 72980
rect 205850 72910 205860 72980
rect 205640 72860 205860 72910
rect 206140 73090 206360 73140
rect 206140 73020 206150 73090
rect 206350 73020 206360 73090
rect 206140 72980 206360 73020
rect 206140 72910 206150 72980
rect 206350 72910 206360 72980
rect 206140 72860 206360 72910
rect 206640 73090 206860 73140
rect 206640 73020 206650 73090
rect 206850 73020 206860 73090
rect 206640 72980 206860 73020
rect 206640 72910 206650 72980
rect 206850 72910 206860 72980
rect 206640 72860 206860 72910
rect 207140 73090 207360 73140
rect 207140 73020 207150 73090
rect 207350 73020 207360 73090
rect 207140 72980 207360 73020
rect 207140 72910 207150 72980
rect 207350 72910 207360 72980
rect 207140 72860 207360 72910
rect 207640 73090 207860 73140
rect 207640 73020 207650 73090
rect 207850 73020 207860 73090
rect 207640 72980 207860 73020
rect 207640 72910 207650 72980
rect 207850 72910 207860 72980
rect 207640 72860 207860 72910
rect 196000 72850 208000 72860
rect 196000 72650 196020 72850
rect 196090 72650 196410 72850
rect 196480 72650 196520 72850
rect 196590 72650 196910 72850
rect 196980 72650 197020 72850
rect 197090 72650 197410 72850
rect 197480 72650 197520 72850
rect 197590 72650 197910 72850
rect 197980 72650 198020 72850
rect 198090 72650 198410 72850
rect 198480 72650 198520 72850
rect 198590 72650 198910 72850
rect 198980 72650 199020 72850
rect 199090 72650 199410 72850
rect 199480 72650 199520 72850
rect 199590 72650 199910 72850
rect 199980 72650 200020 72850
rect 200090 72650 200410 72850
rect 200480 72650 200520 72850
rect 200590 72650 200910 72850
rect 200980 72650 201020 72850
rect 201090 72650 201410 72850
rect 201480 72650 201520 72850
rect 201590 72650 201910 72850
rect 201980 72650 202020 72850
rect 202090 72650 202410 72850
rect 202480 72650 202520 72850
rect 202590 72650 202910 72850
rect 202980 72650 203020 72850
rect 203090 72650 203410 72850
rect 203480 72650 203520 72850
rect 203590 72650 203910 72850
rect 203980 72650 204020 72850
rect 204090 72650 204410 72850
rect 204480 72650 204520 72850
rect 204590 72650 204910 72850
rect 204980 72650 205020 72850
rect 205090 72650 205410 72850
rect 205480 72650 205520 72850
rect 205590 72650 205910 72850
rect 205980 72650 206020 72850
rect 206090 72650 206410 72850
rect 206480 72650 206520 72850
rect 206590 72650 206910 72850
rect 206980 72650 207020 72850
rect 207090 72650 207410 72850
rect 207480 72650 207520 72850
rect 207590 72650 207910 72850
rect 207980 72650 208000 72850
rect 196000 72640 208000 72650
rect 196140 72590 196360 72640
rect 196140 72520 196150 72590
rect 196350 72520 196360 72590
rect 196140 72480 196360 72520
rect 196140 72410 196150 72480
rect 196350 72410 196360 72480
rect 196140 72360 196360 72410
rect 196640 72590 196860 72640
rect 196640 72520 196650 72590
rect 196850 72520 196860 72590
rect 196640 72480 196860 72520
rect 196640 72410 196650 72480
rect 196850 72410 196860 72480
rect 196640 72360 196860 72410
rect 197140 72590 197360 72640
rect 197140 72520 197150 72590
rect 197350 72520 197360 72590
rect 197140 72480 197360 72520
rect 197140 72410 197150 72480
rect 197350 72410 197360 72480
rect 197140 72360 197360 72410
rect 197640 72590 197860 72640
rect 197640 72520 197650 72590
rect 197850 72520 197860 72590
rect 197640 72480 197860 72520
rect 197640 72410 197650 72480
rect 197850 72410 197860 72480
rect 197640 72360 197860 72410
rect 198140 72590 198360 72640
rect 198140 72520 198150 72590
rect 198350 72520 198360 72590
rect 198140 72480 198360 72520
rect 198140 72410 198150 72480
rect 198350 72410 198360 72480
rect 198140 72360 198360 72410
rect 198640 72590 198860 72640
rect 198640 72520 198650 72590
rect 198850 72520 198860 72590
rect 198640 72480 198860 72520
rect 198640 72410 198650 72480
rect 198850 72410 198860 72480
rect 198640 72360 198860 72410
rect 199140 72590 199360 72640
rect 199140 72520 199150 72590
rect 199350 72520 199360 72590
rect 199140 72480 199360 72520
rect 199140 72410 199150 72480
rect 199350 72410 199360 72480
rect 199140 72360 199360 72410
rect 199640 72590 199860 72640
rect 199640 72520 199650 72590
rect 199850 72520 199860 72590
rect 199640 72480 199860 72520
rect 199640 72410 199650 72480
rect 199850 72410 199860 72480
rect 199640 72360 199860 72410
rect 200140 72590 200360 72640
rect 200140 72520 200150 72590
rect 200350 72520 200360 72590
rect 200140 72480 200360 72520
rect 200140 72410 200150 72480
rect 200350 72410 200360 72480
rect 200140 72360 200360 72410
rect 200640 72590 200860 72640
rect 200640 72520 200650 72590
rect 200850 72520 200860 72590
rect 200640 72480 200860 72520
rect 200640 72410 200650 72480
rect 200850 72410 200860 72480
rect 200640 72360 200860 72410
rect 201140 72590 201360 72640
rect 201140 72520 201150 72590
rect 201350 72520 201360 72590
rect 201140 72480 201360 72520
rect 201140 72410 201150 72480
rect 201350 72410 201360 72480
rect 201140 72360 201360 72410
rect 201640 72590 201860 72640
rect 201640 72520 201650 72590
rect 201850 72520 201860 72590
rect 201640 72480 201860 72520
rect 201640 72410 201650 72480
rect 201850 72410 201860 72480
rect 201640 72360 201860 72410
rect 202140 72590 202360 72640
rect 202140 72520 202150 72590
rect 202350 72520 202360 72590
rect 202140 72480 202360 72520
rect 202140 72410 202150 72480
rect 202350 72410 202360 72480
rect 202140 72360 202360 72410
rect 202640 72590 202860 72640
rect 202640 72520 202650 72590
rect 202850 72520 202860 72590
rect 202640 72480 202860 72520
rect 202640 72410 202650 72480
rect 202850 72410 202860 72480
rect 202640 72360 202860 72410
rect 203140 72590 203360 72640
rect 203140 72520 203150 72590
rect 203350 72520 203360 72590
rect 203140 72480 203360 72520
rect 203140 72410 203150 72480
rect 203350 72410 203360 72480
rect 203140 72360 203360 72410
rect 203640 72590 203860 72640
rect 203640 72520 203650 72590
rect 203850 72520 203860 72590
rect 203640 72480 203860 72520
rect 203640 72410 203650 72480
rect 203850 72410 203860 72480
rect 203640 72360 203860 72410
rect 204140 72590 204360 72640
rect 204140 72520 204150 72590
rect 204350 72520 204360 72590
rect 204140 72480 204360 72520
rect 204140 72410 204150 72480
rect 204350 72410 204360 72480
rect 204140 72360 204360 72410
rect 204640 72590 204860 72640
rect 204640 72520 204650 72590
rect 204850 72520 204860 72590
rect 204640 72480 204860 72520
rect 204640 72410 204650 72480
rect 204850 72410 204860 72480
rect 204640 72360 204860 72410
rect 205140 72590 205360 72640
rect 205140 72520 205150 72590
rect 205350 72520 205360 72590
rect 205140 72480 205360 72520
rect 205140 72410 205150 72480
rect 205350 72410 205360 72480
rect 205140 72360 205360 72410
rect 205640 72590 205860 72640
rect 205640 72520 205650 72590
rect 205850 72520 205860 72590
rect 205640 72480 205860 72520
rect 205640 72410 205650 72480
rect 205850 72410 205860 72480
rect 205640 72360 205860 72410
rect 206140 72590 206360 72640
rect 206140 72520 206150 72590
rect 206350 72520 206360 72590
rect 206140 72480 206360 72520
rect 206140 72410 206150 72480
rect 206350 72410 206360 72480
rect 206140 72360 206360 72410
rect 206640 72590 206860 72640
rect 206640 72520 206650 72590
rect 206850 72520 206860 72590
rect 206640 72480 206860 72520
rect 206640 72410 206650 72480
rect 206850 72410 206860 72480
rect 206640 72360 206860 72410
rect 207140 72590 207360 72640
rect 207140 72520 207150 72590
rect 207350 72520 207360 72590
rect 207140 72480 207360 72520
rect 207140 72410 207150 72480
rect 207350 72410 207360 72480
rect 207140 72360 207360 72410
rect 207640 72590 207860 72640
rect 207640 72520 207650 72590
rect 207850 72520 207860 72590
rect 207640 72480 207860 72520
rect 207640 72410 207650 72480
rect 207850 72410 207860 72480
rect 207640 72360 207860 72410
rect 196000 72350 208000 72360
rect 196000 72150 196020 72350
rect 196090 72150 196410 72350
rect 196480 72150 196520 72350
rect 196590 72150 196910 72350
rect 196980 72150 197020 72350
rect 197090 72150 197410 72350
rect 197480 72150 197520 72350
rect 197590 72150 197910 72350
rect 197980 72150 198020 72350
rect 198090 72150 198410 72350
rect 198480 72150 198520 72350
rect 198590 72150 198910 72350
rect 198980 72150 199020 72350
rect 199090 72150 199410 72350
rect 199480 72150 199520 72350
rect 199590 72150 199910 72350
rect 199980 72150 200020 72350
rect 200090 72150 200410 72350
rect 200480 72150 200520 72350
rect 200590 72150 200910 72350
rect 200980 72150 201020 72350
rect 201090 72150 201410 72350
rect 201480 72150 201520 72350
rect 201590 72150 201910 72350
rect 201980 72150 202020 72350
rect 202090 72150 202410 72350
rect 202480 72150 202520 72350
rect 202590 72150 202910 72350
rect 202980 72150 203020 72350
rect 203090 72150 203410 72350
rect 203480 72150 203520 72350
rect 203590 72150 203910 72350
rect 203980 72150 204020 72350
rect 204090 72150 204410 72350
rect 204480 72150 204520 72350
rect 204590 72150 204910 72350
rect 204980 72150 205020 72350
rect 205090 72150 205410 72350
rect 205480 72150 205520 72350
rect 205590 72150 205910 72350
rect 205980 72150 206020 72350
rect 206090 72150 206410 72350
rect 206480 72150 206520 72350
rect 206590 72150 206910 72350
rect 206980 72150 207020 72350
rect 207090 72150 207410 72350
rect 207480 72150 207520 72350
rect 207590 72150 207910 72350
rect 207980 72150 208000 72350
rect 196000 72140 208000 72150
rect 196140 72090 196360 72140
rect 196140 72020 196150 72090
rect 196350 72020 196360 72090
rect 196140 71980 196360 72020
rect 196140 71910 196150 71980
rect 196350 71910 196360 71980
rect 196140 71860 196360 71910
rect 196640 72090 196860 72140
rect 196640 72020 196650 72090
rect 196850 72020 196860 72090
rect 196640 71980 196860 72020
rect 196640 71910 196650 71980
rect 196850 71910 196860 71980
rect 196640 71860 196860 71910
rect 197140 72090 197360 72140
rect 197140 72020 197150 72090
rect 197350 72020 197360 72090
rect 197140 71980 197360 72020
rect 197140 71910 197150 71980
rect 197350 71910 197360 71980
rect 197140 71860 197360 71910
rect 197640 72090 197860 72140
rect 197640 72020 197650 72090
rect 197850 72020 197860 72090
rect 197640 71980 197860 72020
rect 197640 71910 197650 71980
rect 197850 71910 197860 71980
rect 197640 71860 197860 71910
rect 198140 72090 198360 72140
rect 198140 72020 198150 72090
rect 198350 72020 198360 72090
rect 198140 71980 198360 72020
rect 198140 71910 198150 71980
rect 198350 71910 198360 71980
rect 198140 71860 198360 71910
rect 198640 72090 198860 72140
rect 198640 72020 198650 72090
rect 198850 72020 198860 72090
rect 198640 71980 198860 72020
rect 198640 71910 198650 71980
rect 198850 71910 198860 71980
rect 198640 71860 198860 71910
rect 199140 72090 199360 72140
rect 199140 72020 199150 72090
rect 199350 72020 199360 72090
rect 199140 71980 199360 72020
rect 199140 71910 199150 71980
rect 199350 71910 199360 71980
rect 199140 71860 199360 71910
rect 199640 72090 199860 72140
rect 199640 72020 199650 72090
rect 199850 72020 199860 72090
rect 199640 71980 199860 72020
rect 199640 71910 199650 71980
rect 199850 71910 199860 71980
rect 199640 71860 199860 71910
rect 200140 72090 200360 72140
rect 200140 72020 200150 72090
rect 200350 72020 200360 72090
rect 200140 71980 200360 72020
rect 200140 71910 200150 71980
rect 200350 71910 200360 71980
rect 200140 71860 200360 71910
rect 200640 72090 200860 72140
rect 200640 72020 200650 72090
rect 200850 72020 200860 72090
rect 200640 71980 200860 72020
rect 200640 71910 200650 71980
rect 200850 71910 200860 71980
rect 200640 71860 200860 71910
rect 201140 72090 201360 72140
rect 201140 72020 201150 72090
rect 201350 72020 201360 72090
rect 201140 71980 201360 72020
rect 201140 71910 201150 71980
rect 201350 71910 201360 71980
rect 201140 71860 201360 71910
rect 201640 72090 201860 72140
rect 201640 72020 201650 72090
rect 201850 72020 201860 72090
rect 201640 71980 201860 72020
rect 201640 71910 201650 71980
rect 201850 71910 201860 71980
rect 201640 71860 201860 71910
rect 202140 72090 202360 72140
rect 202140 72020 202150 72090
rect 202350 72020 202360 72090
rect 202140 71980 202360 72020
rect 202140 71910 202150 71980
rect 202350 71910 202360 71980
rect 202140 71860 202360 71910
rect 202640 72090 202860 72140
rect 202640 72020 202650 72090
rect 202850 72020 202860 72090
rect 202640 71980 202860 72020
rect 202640 71910 202650 71980
rect 202850 71910 202860 71980
rect 202640 71860 202860 71910
rect 203140 72090 203360 72140
rect 203140 72020 203150 72090
rect 203350 72020 203360 72090
rect 203140 71980 203360 72020
rect 203140 71910 203150 71980
rect 203350 71910 203360 71980
rect 203140 71860 203360 71910
rect 203640 72090 203860 72140
rect 203640 72020 203650 72090
rect 203850 72020 203860 72090
rect 203640 71980 203860 72020
rect 203640 71910 203650 71980
rect 203850 71910 203860 71980
rect 203640 71860 203860 71910
rect 204140 72090 204360 72140
rect 204140 72020 204150 72090
rect 204350 72020 204360 72090
rect 204140 71980 204360 72020
rect 204140 71910 204150 71980
rect 204350 71910 204360 71980
rect 204140 71860 204360 71910
rect 204640 72090 204860 72140
rect 204640 72020 204650 72090
rect 204850 72020 204860 72090
rect 204640 71980 204860 72020
rect 204640 71910 204650 71980
rect 204850 71910 204860 71980
rect 204640 71860 204860 71910
rect 205140 72090 205360 72140
rect 205140 72020 205150 72090
rect 205350 72020 205360 72090
rect 205140 71980 205360 72020
rect 205140 71910 205150 71980
rect 205350 71910 205360 71980
rect 205140 71860 205360 71910
rect 205640 72090 205860 72140
rect 205640 72020 205650 72090
rect 205850 72020 205860 72090
rect 205640 71980 205860 72020
rect 205640 71910 205650 71980
rect 205850 71910 205860 71980
rect 205640 71860 205860 71910
rect 206140 72090 206360 72140
rect 206140 72020 206150 72090
rect 206350 72020 206360 72090
rect 206140 71980 206360 72020
rect 206140 71910 206150 71980
rect 206350 71910 206360 71980
rect 206140 71860 206360 71910
rect 206640 72090 206860 72140
rect 206640 72020 206650 72090
rect 206850 72020 206860 72090
rect 206640 71980 206860 72020
rect 206640 71910 206650 71980
rect 206850 71910 206860 71980
rect 206640 71860 206860 71910
rect 207140 72090 207360 72140
rect 207140 72020 207150 72090
rect 207350 72020 207360 72090
rect 207140 71980 207360 72020
rect 207140 71910 207150 71980
rect 207350 71910 207360 71980
rect 207140 71860 207360 71910
rect 207640 72090 207860 72140
rect 207640 72020 207650 72090
rect 207850 72020 207860 72090
rect 207640 71980 207860 72020
rect 207640 71910 207650 71980
rect 207850 71910 207860 71980
rect 207640 71860 207860 71910
rect 196000 71850 208000 71860
rect 196000 71650 196020 71850
rect 196090 71650 196410 71850
rect 196480 71650 196520 71850
rect 196590 71650 196910 71850
rect 196980 71650 197020 71850
rect 197090 71650 197410 71850
rect 197480 71650 197520 71850
rect 197590 71650 197910 71850
rect 197980 71650 198020 71850
rect 198090 71650 198410 71850
rect 198480 71650 198520 71850
rect 198590 71650 198910 71850
rect 198980 71650 199020 71850
rect 199090 71650 199410 71850
rect 199480 71650 199520 71850
rect 199590 71650 199910 71850
rect 199980 71650 200020 71850
rect 200090 71650 200410 71850
rect 200480 71650 200520 71850
rect 200590 71650 200910 71850
rect 200980 71650 201020 71850
rect 201090 71650 201410 71850
rect 201480 71650 201520 71850
rect 201590 71650 201910 71850
rect 201980 71650 202020 71850
rect 202090 71650 202410 71850
rect 202480 71650 202520 71850
rect 202590 71650 202910 71850
rect 202980 71650 203020 71850
rect 203090 71650 203410 71850
rect 203480 71650 203520 71850
rect 203590 71650 203910 71850
rect 203980 71650 204020 71850
rect 204090 71650 204410 71850
rect 204480 71650 204520 71850
rect 204590 71650 204910 71850
rect 204980 71650 205020 71850
rect 205090 71650 205410 71850
rect 205480 71650 205520 71850
rect 205590 71650 205910 71850
rect 205980 71650 206020 71850
rect 206090 71650 206410 71850
rect 206480 71650 206520 71850
rect 206590 71650 206910 71850
rect 206980 71650 207020 71850
rect 207090 71650 207410 71850
rect 207480 71650 207520 71850
rect 207590 71650 207910 71850
rect 207980 71650 208000 71850
rect 196000 71640 208000 71650
rect 196140 71590 196360 71640
rect 196140 71520 196150 71590
rect 196350 71520 196360 71590
rect 196140 71480 196360 71520
rect 196140 71410 196150 71480
rect 196350 71410 196360 71480
rect 196140 71360 196360 71410
rect 196640 71590 196860 71640
rect 196640 71520 196650 71590
rect 196850 71520 196860 71590
rect 196640 71480 196860 71520
rect 196640 71410 196650 71480
rect 196850 71410 196860 71480
rect 196640 71360 196860 71410
rect 197140 71590 197360 71640
rect 197140 71520 197150 71590
rect 197350 71520 197360 71590
rect 197140 71480 197360 71520
rect 197140 71410 197150 71480
rect 197350 71410 197360 71480
rect 197140 71360 197360 71410
rect 197640 71590 197860 71640
rect 197640 71520 197650 71590
rect 197850 71520 197860 71590
rect 197640 71480 197860 71520
rect 197640 71410 197650 71480
rect 197850 71410 197860 71480
rect 197640 71360 197860 71410
rect 198140 71590 198360 71640
rect 198140 71520 198150 71590
rect 198350 71520 198360 71590
rect 198140 71480 198360 71520
rect 198140 71410 198150 71480
rect 198350 71410 198360 71480
rect 198140 71360 198360 71410
rect 198640 71590 198860 71640
rect 198640 71520 198650 71590
rect 198850 71520 198860 71590
rect 198640 71480 198860 71520
rect 198640 71410 198650 71480
rect 198850 71410 198860 71480
rect 198640 71360 198860 71410
rect 199140 71590 199360 71640
rect 199140 71520 199150 71590
rect 199350 71520 199360 71590
rect 199140 71480 199360 71520
rect 199140 71410 199150 71480
rect 199350 71410 199360 71480
rect 199140 71360 199360 71410
rect 199640 71590 199860 71640
rect 199640 71520 199650 71590
rect 199850 71520 199860 71590
rect 199640 71480 199860 71520
rect 199640 71410 199650 71480
rect 199850 71410 199860 71480
rect 199640 71360 199860 71410
rect 200140 71590 200360 71640
rect 200140 71520 200150 71590
rect 200350 71520 200360 71590
rect 200140 71480 200360 71520
rect 200140 71410 200150 71480
rect 200350 71410 200360 71480
rect 200140 71360 200360 71410
rect 200640 71590 200860 71640
rect 200640 71520 200650 71590
rect 200850 71520 200860 71590
rect 200640 71480 200860 71520
rect 200640 71410 200650 71480
rect 200850 71410 200860 71480
rect 200640 71360 200860 71410
rect 201140 71590 201360 71640
rect 201140 71520 201150 71590
rect 201350 71520 201360 71590
rect 201140 71480 201360 71520
rect 201140 71410 201150 71480
rect 201350 71410 201360 71480
rect 201140 71360 201360 71410
rect 201640 71590 201860 71640
rect 201640 71520 201650 71590
rect 201850 71520 201860 71590
rect 201640 71480 201860 71520
rect 201640 71410 201650 71480
rect 201850 71410 201860 71480
rect 201640 71360 201860 71410
rect 202140 71590 202360 71640
rect 202140 71520 202150 71590
rect 202350 71520 202360 71590
rect 202140 71480 202360 71520
rect 202140 71410 202150 71480
rect 202350 71410 202360 71480
rect 202140 71360 202360 71410
rect 202640 71590 202860 71640
rect 202640 71520 202650 71590
rect 202850 71520 202860 71590
rect 202640 71480 202860 71520
rect 202640 71410 202650 71480
rect 202850 71410 202860 71480
rect 202640 71360 202860 71410
rect 203140 71590 203360 71640
rect 203140 71520 203150 71590
rect 203350 71520 203360 71590
rect 203140 71480 203360 71520
rect 203140 71410 203150 71480
rect 203350 71410 203360 71480
rect 203140 71360 203360 71410
rect 203640 71590 203860 71640
rect 203640 71520 203650 71590
rect 203850 71520 203860 71590
rect 203640 71480 203860 71520
rect 203640 71410 203650 71480
rect 203850 71410 203860 71480
rect 203640 71360 203860 71410
rect 204140 71590 204360 71640
rect 204140 71520 204150 71590
rect 204350 71520 204360 71590
rect 204140 71480 204360 71520
rect 204140 71410 204150 71480
rect 204350 71410 204360 71480
rect 204140 71360 204360 71410
rect 204640 71590 204860 71640
rect 204640 71520 204650 71590
rect 204850 71520 204860 71590
rect 204640 71480 204860 71520
rect 204640 71410 204650 71480
rect 204850 71410 204860 71480
rect 204640 71360 204860 71410
rect 205140 71590 205360 71640
rect 205140 71520 205150 71590
rect 205350 71520 205360 71590
rect 205140 71480 205360 71520
rect 205140 71410 205150 71480
rect 205350 71410 205360 71480
rect 205140 71360 205360 71410
rect 205640 71590 205860 71640
rect 205640 71520 205650 71590
rect 205850 71520 205860 71590
rect 205640 71480 205860 71520
rect 205640 71410 205650 71480
rect 205850 71410 205860 71480
rect 205640 71360 205860 71410
rect 206140 71590 206360 71640
rect 206140 71520 206150 71590
rect 206350 71520 206360 71590
rect 206140 71480 206360 71520
rect 206140 71410 206150 71480
rect 206350 71410 206360 71480
rect 206140 71360 206360 71410
rect 206640 71590 206860 71640
rect 206640 71520 206650 71590
rect 206850 71520 206860 71590
rect 206640 71480 206860 71520
rect 206640 71410 206650 71480
rect 206850 71410 206860 71480
rect 206640 71360 206860 71410
rect 207140 71590 207360 71640
rect 207140 71520 207150 71590
rect 207350 71520 207360 71590
rect 207140 71480 207360 71520
rect 207140 71410 207150 71480
rect 207350 71410 207360 71480
rect 207140 71360 207360 71410
rect 207640 71590 207860 71640
rect 207640 71520 207650 71590
rect 207850 71520 207860 71590
rect 207640 71480 207860 71520
rect 207640 71410 207650 71480
rect 207850 71410 207860 71480
rect 207640 71360 207860 71410
rect 196000 71350 208000 71360
rect 196000 71150 196020 71350
rect 196090 71150 196410 71350
rect 196480 71150 196520 71350
rect 196590 71150 196910 71350
rect 196980 71150 197020 71350
rect 197090 71150 197410 71350
rect 197480 71150 197520 71350
rect 197590 71150 197910 71350
rect 197980 71150 198020 71350
rect 198090 71150 198410 71350
rect 198480 71150 198520 71350
rect 198590 71150 198910 71350
rect 198980 71150 199020 71350
rect 199090 71150 199410 71350
rect 199480 71150 199520 71350
rect 199590 71150 199910 71350
rect 199980 71150 200020 71350
rect 200090 71150 200410 71350
rect 200480 71150 200520 71350
rect 200590 71150 200910 71350
rect 200980 71150 201020 71350
rect 201090 71150 201410 71350
rect 201480 71150 201520 71350
rect 201590 71150 201910 71350
rect 201980 71150 202020 71350
rect 202090 71150 202410 71350
rect 202480 71150 202520 71350
rect 202590 71150 202910 71350
rect 202980 71150 203020 71350
rect 203090 71150 203410 71350
rect 203480 71150 203520 71350
rect 203590 71150 203910 71350
rect 203980 71150 204020 71350
rect 204090 71150 204410 71350
rect 204480 71150 204520 71350
rect 204590 71150 204910 71350
rect 204980 71150 205020 71350
rect 205090 71150 205410 71350
rect 205480 71150 205520 71350
rect 205590 71150 205910 71350
rect 205980 71150 206020 71350
rect 206090 71150 206410 71350
rect 206480 71150 206520 71350
rect 206590 71150 206910 71350
rect 206980 71150 207020 71350
rect 207090 71150 207410 71350
rect 207480 71150 207520 71350
rect 207590 71150 207910 71350
rect 207980 71150 208000 71350
rect 196000 71140 208000 71150
rect 196140 71090 196360 71140
rect 196140 71020 196150 71090
rect 196350 71020 196360 71090
rect 196140 70980 196360 71020
rect 196140 70910 196150 70980
rect 196350 70910 196360 70980
rect 196140 70860 196360 70910
rect 196640 71090 196860 71140
rect 196640 71020 196650 71090
rect 196850 71020 196860 71090
rect 196640 70980 196860 71020
rect 196640 70910 196650 70980
rect 196850 70910 196860 70980
rect 196640 70860 196860 70910
rect 197140 71090 197360 71140
rect 197140 71020 197150 71090
rect 197350 71020 197360 71090
rect 197140 70980 197360 71020
rect 197140 70910 197150 70980
rect 197350 70910 197360 70980
rect 197140 70860 197360 70910
rect 197640 71090 197860 71140
rect 197640 71020 197650 71090
rect 197850 71020 197860 71090
rect 197640 70980 197860 71020
rect 197640 70910 197650 70980
rect 197850 70910 197860 70980
rect 197640 70860 197860 70910
rect 198140 71090 198360 71140
rect 198140 71020 198150 71090
rect 198350 71020 198360 71090
rect 198140 70980 198360 71020
rect 198140 70910 198150 70980
rect 198350 70910 198360 70980
rect 198140 70860 198360 70910
rect 198640 71090 198860 71140
rect 198640 71020 198650 71090
rect 198850 71020 198860 71090
rect 198640 70980 198860 71020
rect 198640 70910 198650 70980
rect 198850 70910 198860 70980
rect 198640 70860 198860 70910
rect 199140 71090 199360 71140
rect 199140 71020 199150 71090
rect 199350 71020 199360 71090
rect 199140 70980 199360 71020
rect 199140 70910 199150 70980
rect 199350 70910 199360 70980
rect 199140 70860 199360 70910
rect 199640 71090 199860 71140
rect 199640 71020 199650 71090
rect 199850 71020 199860 71090
rect 199640 70980 199860 71020
rect 199640 70910 199650 70980
rect 199850 70910 199860 70980
rect 199640 70860 199860 70910
rect 200140 71090 200360 71140
rect 200140 71020 200150 71090
rect 200350 71020 200360 71090
rect 200140 70980 200360 71020
rect 200140 70910 200150 70980
rect 200350 70910 200360 70980
rect 200140 70860 200360 70910
rect 200640 71090 200860 71140
rect 200640 71020 200650 71090
rect 200850 71020 200860 71090
rect 200640 70980 200860 71020
rect 200640 70910 200650 70980
rect 200850 70910 200860 70980
rect 200640 70860 200860 70910
rect 201140 71090 201360 71140
rect 201140 71020 201150 71090
rect 201350 71020 201360 71090
rect 201140 70980 201360 71020
rect 201140 70910 201150 70980
rect 201350 70910 201360 70980
rect 201140 70860 201360 70910
rect 201640 71090 201860 71140
rect 201640 71020 201650 71090
rect 201850 71020 201860 71090
rect 201640 70980 201860 71020
rect 201640 70910 201650 70980
rect 201850 70910 201860 70980
rect 201640 70860 201860 70910
rect 202140 71090 202360 71140
rect 202140 71020 202150 71090
rect 202350 71020 202360 71090
rect 202140 70980 202360 71020
rect 202140 70910 202150 70980
rect 202350 70910 202360 70980
rect 202140 70860 202360 70910
rect 202640 71090 202860 71140
rect 202640 71020 202650 71090
rect 202850 71020 202860 71090
rect 202640 70980 202860 71020
rect 202640 70910 202650 70980
rect 202850 70910 202860 70980
rect 202640 70860 202860 70910
rect 203140 71090 203360 71140
rect 203140 71020 203150 71090
rect 203350 71020 203360 71090
rect 203140 70980 203360 71020
rect 203140 70910 203150 70980
rect 203350 70910 203360 70980
rect 203140 70860 203360 70910
rect 203640 71090 203860 71140
rect 203640 71020 203650 71090
rect 203850 71020 203860 71090
rect 203640 70980 203860 71020
rect 203640 70910 203650 70980
rect 203850 70910 203860 70980
rect 203640 70860 203860 70910
rect 204140 71090 204360 71140
rect 204140 71020 204150 71090
rect 204350 71020 204360 71090
rect 204140 70980 204360 71020
rect 204140 70910 204150 70980
rect 204350 70910 204360 70980
rect 204140 70860 204360 70910
rect 204640 71090 204860 71140
rect 204640 71020 204650 71090
rect 204850 71020 204860 71090
rect 204640 70980 204860 71020
rect 204640 70910 204650 70980
rect 204850 70910 204860 70980
rect 204640 70860 204860 70910
rect 205140 71090 205360 71140
rect 205140 71020 205150 71090
rect 205350 71020 205360 71090
rect 205140 70980 205360 71020
rect 205140 70910 205150 70980
rect 205350 70910 205360 70980
rect 205140 70860 205360 70910
rect 205640 71090 205860 71140
rect 205640 71020 205650 71090
rect 205850 71020 205860 71090
rect 205640 70980 205860 71020
rect 205640 70910 205650 70980
rect 205850 70910 205860 70980
rect 205640 70860 205860 70910
rect 206140 71090 206360 71140
rect 206140 71020 206150 71090
rect 206350 71020 206360 71090
rect 206140 70980 206360 71020
rect 206140 70910 206150 70980
rect 206350 70910 206360 70980
rect 206140 70860 206360 70910
rect 206640 71090 206860 71140
rect 206640 71020 206650 71090
rect 206850 71020 206860 71090
rect 206640 70980 206860 71020
rect 206640 70910 206650 70980
rect 206850 70910 206860 70980
rect 206640 70860 206860 70910
rect 207140 71090 207360 71140
rect 207140 71020 207150 71090
rect 207350 71020 207360 71090
rect 207140 70980 207360 71020
rect 207140 70910 207150 70980
rect 207350 70910 207360 70980
rect 207140 70860 207360 70910
rect 207640 71090 207860 71140
rect 207640 71020 207650 71090
rect 207850 71020 207860 71090
rect 207640 70980 207860 71020
rect 207640 70910 207650 70980
rect 207850 70910 207860 70980
rect 207640 70860 207860 70910
rect 196000 70850 208000 70860
rect 196000 70650 196020 70850
rect 196090 70650 196410 70850
rect 196480 70650 196520 70850
rect 196590 70650 196910 70850
rect 196980 70650 197020 70850
rect 197090 70650 197410 70850
rect 197480 70650 197520 70850
rect 197590 70650 197910 70850
rect 197980 70650 198020 70850
rect 198090 70650 198410 70850
rect 198480 70650 198520 70850
rect 198590 70650 198910 70850
rect 198980 70650 199020 70850
rect 199090 70650 199410 70850
rect 199480 70650 199520 70850
rect 199590 70650 199910 70850
rect 199980 70650 200020 70850
rect 200090 70650 200410 70850
rect 200480 70650 200520 70850
rect 200590 70650 200910 70850
rect 200980 70650 201020 70850
rect 201090 70650 201410 70850
rect 201480 70650 201520 70850
rect 201590 70650 201910 70850
rect 201980 70650 202020 70850
rect 202090 70650 202410 70850
rect 202480 70650 202520 70850
rect 202590 70650 202910 70850
rect 202980 70650 203020 70850
rect 203090 70650 203410 70850
rect 203480 70650 203520 70850
rect 203590 70650 203910 70850
rect 203980 70650 204020 70850
rect 204090 70650 204410 70850
rect 204480 70650 204520 70850
rect 204590 70650 204910 70850
rect 204980 70650 205020 70850
rect 205090 70650 205410 70850
rect 205480 70650 205520 70850
rect 205590 70650 205910 70850
rect 205980 70650 206020 70850
rect 206090 70650 206410 70850
rect 206480 70650 206520 70850
rect 206590 70650 206910 70850
rect 206980 70650 207020 70850
rect 207090 70650 207410 70850
rect 207480 70650 207520 70850
rect 207590 70650 207910 70850
rect 207980 70650 208000 70850
rect 196000 70640 208000 70650
rect 196140 70590 196360 70640
rect 196140 70520 196150 70590
rect 196350 70520 196360 70590
rect 196140 70480 196360 70520
rect 196140 70410 196150 70480
rect 196350 70410 196360 70480
rect 196140 70360 196360 70410
rect 196640 70590 196860 70640
rect 196640 70520 196650 70590
rect 196850 70520 196860 70590
rect 196640 70480 196860 70520
rect 196640 70410 196650 70480
rect 196850 70410 196860 70480
rect 196640 70360 196860 70410
rect 197140 70590 197360 70640
rect 197140 70520 197150 70590
rect 197350 70520 197360 70590
rect 197140 70480 197360 70520
rect 197140 70410 197150 70480
rect 197350 70410 197360 70480
rect 197140 70360 197360 70410
rect 197640 70590 197860 70640
rect 197640 70520 197650 70590
rect 197850 70520 197860 70590
rect 197640 70480 197860 70520
rect 197640 70410 197650 70480
rect 197850 70410 197860 70480
rect 197640 70360 197860 70410
rect 198140 70590 198360 70640
rect 198140 70520 198150 70590
rect 198350 70520 198360 70590
rect 198140 70480 198360 70520
rect 198140 70410 198150 70480
rect 198350 70410 198360 70480
rect 198140 70360 198360 70410
rect 198640 70590 198860 70640
rect 198640 70520 198650 70590
rect 198850 70520 198860 70590
rect 198640 70480 198860 70520
rect 198640 70410 198650 70480
rect 198850 70410 198860 70480
rect 198640 70360 198860 70410
rect 199140 70590 199360 70640
rect 199140 70520 199150 70590
rect 199350 70520 199360 70590
rect 199140 70480 199360 70520
rect 199140 70410 199150 70480
rect 199350 70410 199360 70480
rect 199140 70360 199360 70410
rect 199640 70590 199860 70640
rect 199640 70520 199650 70590
rect 199850 70520 199860 70590
rect 199640 70480 199860 70520
rect 199640 70410 199650 70480
rect 199850 70410 199860 70480
rect 199640 70360 199860 70410
rect 200140 70590 200360 70640
rect 200140 70520 200150 70590
rect 200350 70520 200360 70590
rect 200140 70480 200360 70520
rect 200140 70410 200150 70480
rect 200350 70410 200360 70480
rect 200140 70360 200360 70410
rect 200640 70590 200860 70640
rect 200640 70520 200650 70590
rect 200850 70520 200860 70590
rect 200640 70480 200860 70520
rect 200640 70410 200650 70480
rect 200850 70410 200860 70480
rect 200640 70360 200860 70410
rect 201140 70590 201360 70640
rect 201140 70520 201150 70590
rect 201350 70520 201360 70590
rect 201140 70480 201360 70520
rect 201140 70410 201150 70480
rect 201350 70410 201360 70480
rect 201140 70360 201360 70410
rect 201640 70590 201860 70640
rect 201640 70520 201650 70590
rect 201850 70520 201860 70590
rect 201640 70480 201860 70520
rect 201640 70410 201650 70480
rect 201850 70410 201860 70480
rect 201640 70360 201860 70410
rect 202140 70590 202360 70640
rect 202140 70520 202150 70590
rect 202350 70520 202360 70590
rect 202140 70480 202360 70520
rect 202140 70410 202150 70480
rect 202350 70410 202360 70480
rect 202140 70360 202360 70410
rect 202640 70590 202860 70640
rect 202640 70520 202650 70590
rect 202850 70520 202860 70590
rect 202640 70480 202860 70520
rect 202640 70410 202650 70480
rect 202850 70410 202860 70480
rect 202640 70360 202860 70410
rect 203140 70590 203360 70640
rect 203140 70520 203150 70590
rect 203350 70520 203360 70590
rect 203140 70480 203360 70520
rect 203140 70410 203150 70480
rect 203350 70410 203360 70480
rect 203140 70360 203360 70410
rect 203640 70590 203860 70640
rect 203640 70520 203650 70590
rect 203850 70520 203860 70590
rect 203640 70480 203860 70520
rect 203640 70410 203650 70480
rect 203850 70410 203860 70480
rect 203640 70360 203860 70410
rect 204140 70590 204360 70640
rect 204140 70520 204150 70590
rect 204350 70520 204360 70590
rect 204140 70480 204360 70520
rect 204140 70410 204150 70480
rect 204350 70410 204360 70480
rect 204140 70360 204360 70410
rect 204640 70590 204860 70640
rect 204640 70520 204650 70590
rect 204850 70520 204860 70590
rect 204640 70480 204860 70520
rect 204640 70410 204650 70480
rect 204850 70410 204860 70480
rect 204640 70360 204860 70410
rect 205140 70590 205360 70640
rect 205140 70520 205150 70590
rect 205350 70520 205360 70590
rect 205140 70480 205360 70520
rect 205140 70410 205150 70480
rect 205350 70410 205360 70480
rect 205140 70360 205360 70410
rect 205640 70590 205860 70640
rect 205640 70520 205650 70590
rect 205850 70520 205860 70590
rect 205640 70480 205860 70520
rect 205640 70410 205650 70480
rect 205850 70410 205860 70480
rect 205640 70360 205860 70410
rect 206140 70590 206360 70640
rect 206140 70520 206150 70590
rect 206350 70520 206360 70590
rect 206140 70480 206360 70520
rect 206140 70410 206150 70480
rect 206350 70410 206360 70480
rect 206140 70360 206360 70410
rect 206640 70590 206860 70640
rect 206640 70520 206650 70590
rect 206850 70520 206860 70590
rect 206640 70480 206860 70520
rect 206640 70410 206650 70480
rect 206850 70410 206860 70480
rect 206640 70360 206860 70410
rect 207140 70590 207360 70640
rect 207140 70520 207150 70590
rect 207350 70520 207360 70590
rect 207140 70480 207360 70520
rect 207140 70410 207150 70480
rect 207350 70410 207360 70480
rect 207140 70360 207360 70410
rect 207640 70590 207860 70640
rect 207640 70520 207650 70590
rect 207850 70520 207860 70590
rect 207640 70480 207860 70520
rect 207640 70410 207650 70480
rect 207850 70410 207860 70480
rect 207640 70360 207860 70410
rect 196000 70350 208000 70360
rect 196000 70150 196020 70350
rect 196090 70150 196410 70350
rect 196480 70150 196520 70350
rect 196590 70150 196910 70350
rect 196980 70150 197020 70350
rect 197090 70150 197410 70350
rect 197480 70150 197520 70350
rect 197590 70150 197910 70350
rect 197980 70150 198020 70350
rect 198090 70150 198410 70350
rect 198480 70150 198520 70350
rect 198590 70150 198910 70350
rect 198980 70150 199020 70350
rect 199090 70150 199410 70350
rect 199480 70150 199520 70350
rect 199590 70150 199910 70350
rect 199980 70150 200020 70350
rect 200090 70150 200410 70350
rect 200480 70150 200520 70350
rect 200590 70150 200910 70350
rect 200980 70150 201020 70350
rect 201090 70150 201410 70350
rect 201480 70150 201520 70350
rect 201590 70150 201910 70350
rect 201980 70150 202020 70350
rect 202090 70150 202410 70350
rect 202480 70150 202520 70350
rect 202590 70150 202910 70350
rect 202980 70150 203020 70350
rect 203090 70150 203410 70350
rect 203480 70150 203520 70350
rect 203590 70150 203910 70350
rect 203980 70150 204020 70350
rect 204090 70150 204410 70350
rect 204480 70150 204520 70350
rect 204590 70150 204910 70350
rect 204980 70150 205020 70350
rect 205090 70150 205410 70350
rect 205480 70150 205520 70350
rect 205590 70150 205910 70350
rect 205980 70150 206020 70350
rect 206090 70150 206410 70350
rect 206480 70150 206520 70350
rect 206590 70150 206910 70350
rect 206980 70150 207020 70350
rect 207090 70150 207410 70350
rect 207480 70150 207520 70350
rect 207590 70150 207910 70350
rect 207980 70150 208000 70350
rect 196000 70140 208000 70150
rect 196140 70090 196360 70140
rect 196140 70020 196150 70090
rect 196350 70020 196360 70090
rect 196140 69980 196360 70020
rect 196140 69910 196150 69980
rect 196350 69910 196360 69980
rect 196140 69860 196360 69910
rect 196640 70090 196860 70140
rect 196640 70020 196650 70090
rect 196850 70020 196860 70090
rect 196640 69980 196860 70020
rect 196640 69910 196650 69980
rect 196850 69910 196860 69980
rect 196640 69860 196860 69910
rect 197140 70090 197360 70140
rect 197140 70020 197150 70090
rect 197350 70020 197360 70090
rect 197140 69980 197360 70020
rect 197140 69910 197150 69980
rect 197350 69910 197360 69980
rect 197140 69860 197360 69910
rect 197640 70090 197860 70140
rect 197640 70020 197650 70090
rect 197850 70020 197860 70090
rect 197640 69980 197860 70020
rect 197640 69910 197650 69980
rect 197850 69910 197860 69980
rect 197640 69860 197860 69910
rect 198140 70090 198360 70140
rect 198140 70020 198150 70090
rect 198350 70020 198360 70090
rect 198140 69980 198360 70020
rect 198140 69910 198150 69980
rect 198350 69910 198360 69980
rect 198140 69860 198360 69910
rect 198640 70090 198860 70140
rect 198640 70020 198650 70090
rect 198850 70020 198860 70090
rect 198640 69980 198860 70020
rect 198640 69910 198650 69980
rect 198850 69910 198860 69980
rect 198640 69860 198860 69910
rect 199140 70090 199360 70140
rect 199140 70020 199150 70090
rect 199350 70020 199360 70090
rect 199140 69980 199360 70020
rect 199140 69910 199150 69980
rect 199350 69910 199360 69980
rect 199140 69860 199360 69910
rect 199640 70090 199860 70140
rect 199640 70020 199650 70090
rect 199850 70020 199860 70090
rect 199640 69980 199860 70020
rect 199640 69910 199650 69980
rect 199850 69910 199860 69980
rect 199640 69860 199860 69910
rect 200140 70090 200360 70140
rect 200140 70020 200150 70090
rect 200350 70020 200360 70090
rect 200140 69980 200360 70020
rect 200140 69910 200150 69980
rect 200350 69910 200360 69980
rect 200140 69860 200360 69910
rect 200640 70090 200860 70140
rect 200640 70020 200650 70090
rect 200850 70020 200860 70090
rect 200640 69980 200860 70020
rect 200640 69910 200650 69980
rect 200850 69910 200860 69980
rect 200640 69860 200860 69910
rect 201140 70090 201360 70140
rect 201140 70020 201150 70090
rect 201350 70020 201360 70090
rect 201140 69980 201360 70020
rect 201140 69910 201150 69980
rect 201350 69910 201360 69980
rect 201140 69860 201360 69910
rect 201640 70090 201860 70140
rect 201640 70020 201650 70090
rect 201850 70020 201860 70090
rect 201640 69980 201860 70020
rect 201640 69910 201650 69980
rect 201850 69910 201860 69980
rect 201640 69860 201860 69910
rect 202140 70090 202360 70140
rect 202140 70020 202150 70090
rect 202350 70020 202360 70090
rect 202140 69980 202360 70020
rect 202140 69910 202150 69980
rect 202350 69910 202360 69980
rect 202140 69860 202360 69910
rect 202640 70090 202860 70140
rect 202640 70020 202650 70090
rect 202850 70020 202860 70090
rect 202640 69980 202860 70020
rect 202640 69910 202650 69980
rect 202850 69910 202860 69980
rect 202640 69860 202860 69910
rect 203140 70090 203360 70140
rect 203140 70020 203150 70090
rect 203350 70020 203360 70090
rect 203140 69980 203360 70020
rect 203140 69910 203150 69980
rect 203350 69910 203360 69980
rect 203140 69860 203360 69910
rect 203640 70090 203860 70140
rect 203640 70020 203650 70090
rect 203850 70020 203860 70090
rect 203640 69980 203860 70020
rect 203640 69910 203650 69980
rect 203850 69910 203860 69980
rect 203640 69860 203860 69910
rect 204140 70090 204360 70140
rect 204140 70020 204150 70090
rect 204350 70020 204360 70090
rect 204140 69980 204360 70020
rect 204140 69910 204150 69980
rect 204350 69910 204360 69980
rect 204140 69860 204360 69910
rect 204640 70090 204860 70140
rect 204640 70020 204650 70090
rect 204850 70020 204860 70090
rect 204640 69980 204860 70020
rect 204640 69910 204650 69980
rect 204850 69910 204860 69980
rect 204640 69860 204860 69910
rect 205140 70090 205360 70140
rect 205140 70020 205150 70090
rect 205350 70020 205360 70090
rect 205140 69980 205360 70020
rect 205140 69910 205150 69980
rect 205350 69910 205360 69980
rect 205140 69860 205360 69910
rect 205640 70090 205860 70140
rect 205640 70020 205650 70090
rect 205850 70020 205860 70090
rect 205640 69980 205860 70020
rect 205640 69910 205650 69980
rect 205850 69910 205860 69980
rect 205640 69860 205860 69910
rect 206140 70090 206360 70140
rect 206140 70020 206150 70090
rect 206350 70020 206360 70090
rect 206140 69980 206360 70020
rect 206140 69910 206150 69980
rect 206350 69910 206360 69980
rect 206140 69860 206360 69910
rect 206640 70090 206860 70140
rect 206640 70020 206650 70090
rect 206850 70020 206860 70090
rect 206640 69980 206860 70020
rect 206640 69910 206650 69980
rect 206850 69910 206860 69980
rect 206640 69860 206860 69910
rect 207140 70090 207360 70140
rect 207140 70020 207150 70090
rect 207350 70020 207360 70090
rect 207140 69980 207360 70020
rect 207140 69910 207150 69980
rect 207350 69910 207360 69980
rect 207140 69860 207360 69910
rect 207640 70090 207860 70140
rect 207640 70020 207650 70090
rect 207850 70020 207860 70090
rect 207640 69980 207860 70020
rect 207640 69910 207650 69980
rect 207850 69910 207860 69980
rect 207640 69860 207860 69910
rect 196000 69850 208000 69860
rect 196000 69650 196020 69850
rect 196090 69650 196410 69850
rect 196480 69650 196520 69850
rect 196590 69650 196910 69850
rect 196980 69650 197020 69850
rect 197090 69650 197410 69850
rect 197480 69650 197520 69850
rect 197590 69650 197910 69850
rect 197980 69650 198020 69850
rect 198090 69650 198410 69850
rect 198480 69650 198520 69850
rect 198590 69650 198910 69850
rect 198980 69650 199020 69850
rect 199090 69650 199410 69850
rect 199480 69650 199520 69850
rect 199590 69650 199910 69850
rect 199980 69650 200020 69850
rect 200090 69650 200410 69850
rect 200480 69650 200520 69850
rect 200590 69650 200910 69850
rect 200980 69650 201020 69850
rect 201090 69650 201410 69850
rect 201480 69650 201520 69850
rect 201590 69650 201910 69850
rect 201980 69650 202020 69850
rect 202090 69650 202410 69850
rect 202480 69650 202520 69850
rect 202590 69650 202910 69850
rect 202980 69650 203020 69850
rect 203090 69650 203410 69850
rect 203480 69650 203520 69850
rect 203590 69650 203910 69850
rect 203980 69650 204020 69850
rect 204090 69650 204410 69850
rect 204480 69650 204520 69850
rect 204590 69650 204910 69850
rect 204980 69650 205020 69850
rect 205090 69650 205410 69850
rect 205480 69650 205520 69850
rect 205590 69650 205910 69850
rect 205980 69650 206020 69850
rect 206090 69650 206410 69850
rect 206480 69650 206520 69850
rect 206590 69650 206910 69850
rect 206980 69650 207020 69850
rect 207090 69650 207410 69850
rect 207480 69650 207520 69850
rect 207590 69650 207910 69850
rect 207980 69650 208000 69850
rect 196000 69640 208000 69650
rect 196140 69590 196360 69640
rect 196140 69520 196150 69590
rect 196350 69520 196360 69590
rect 196140 69480 196360 69520
rect 196140 69410 196150 69480
rect 196350 69410 196360 69480
rect 196140 69360 196360 69410
rect 196640 69590 196860 69640
rect 196640 69520 196650 69590
rect 196850 69520 196860 69590
rect 196640 69480 196860 69520
rect 196640 69410 196650 69480
rect 196850 69410 196860 69480
rect 196640 69360 196860 69410
rect 197140 69590 197360 69640
rect 197140 69520 197150 69590
rect 197350 69520 197360 69590
rect 197140 69480 197360 69520
rect 197140 69410 197150 69480
rect 197350 69410 197360 69480
rect 197140 69360 197360 69410
rect 197640 69590 197860 69640
rect 197640 69520 197650 69590
rect 197850 69520 197860 69590
rect 197640 69480 197860 69520
rect 197640 69410 197650 69480
rect 197850 69410 197860 69480
rect 197640 69360 197860 69410
rect 198140 69590 198360 69640
rect 198140 69520 198150 69590
rect 198350 69520 198360 69590
rect 198140 69480 198360 69520
rect 198140 69410 198150 69480
rect 198350 69410 198360 69480
rect 198140 69360 198360 69410
rect 198640 69590 198860 69640
rect 198640 69520 198650 69590
rect 198850 69520 198860 69590
rect 198640 69480 198860 69520
rect 198640 69410 198650 69480
rect 198850 69410 198860 69480
rect 198640 69360 198860 69410
rect 199140 69590 199360 69640
rect 199140 69520 199150 69590
rect 199350 69520 199360 69590
rect 199140 69480 199360 69520
rect 199140 69410 199150 69480
rect 199350 69410 199360 69480
rect 199140 69360 199360 69410
rect 199640 69590 199860 69640
rect 199640 69520 199650 69590
rect 199850 69520 199860 69590
rect 199640 69480 199860 69520
rect 199640 69410 199650 69480
rect 199850 69410 199860 69480
rect 199640 69360 199860 69410
rect 200140 69590 200360 69640
rect 200140 69520 200150 69590
rect 200350 69520 200360 69590
rect 200140 69480 200360 69520
rect 200140 69410 200150 69480
rect 200350 69410 200360 69480
rect 200140 69360 200360 69410
rect 200640 69590 200860 69640
rect 200640 69520 200650 69590
rect 200850 69520 200860 69590
rect 200640 69480 200860 69520
rect 200640 69410 200650 69480
rect 200850 69410 200860 69480
rect 200640 69360 200860 69410
rect 201140 69590 201360 69640
rect 201140 69520 201150 69590
rect 201350 69520 201360 69590
rect 201140 69480 201360 69520
rect 201140 69410 201150 69480
rect 201350 69410 201360 69480
rect 201140 69360 201360 69410
rect 201640 69590 201860 69640
rect 201640 69520 201650 69590
rect 201850 69520 201860 69590
rect 201640 69480 201860 69520
rect 201640 69410 201650 69480
rect 201850 69410 201860 69480
rect 201640 69360 201860 69410
rect 202140 69590 202360 69640
rect 202140 69520 202150 69590
rect 202350 69520 202360 69590
rect 202140 69480 202360 69520
rect 202140 69410 202150 69480
rect 202350 69410 202360 69480
rect 202140 69360 202360 69410
rect 202640 69590 202860 69640
rect 202640 69520 202650 69590
rect 202850 69520 202860 69590
rect 202640 69480 202860 69520
rect 202640 69410 202650 69480
rect 202850 69410 202860 69480
rect 202640 69360 202860 69410
rect 203140 69590 203360 69640
rect 203140 69520 203150 69590
rect 203350 69520 203360 69590
rect 203140 69480 203360 69520
rect 203140 69410 203150 69480
rect 203350 69410 203360 69480
rect 203140 69360 203360 69410
rect 203640 69590 203860 69640
rect 203640 69520 203650 69590
rect 203850 69520 203860 69590
rect 203640 69480 203860 69520
rect 203640 69410 203650 69480
rect 203850 69410 203860 69480
rect 203640 69360 203860 69410
rect 204140 69590 204360 69640
rect 204140 69520 204150 69590
rect 204350 69520 204360 69590
rect 204140 69480 204360 69520
rect 204140 69410 204150 69480
rect 204350 69410 204360 69480
rect 204140 69360 204360 69410
rect 204640 69590 204860 69640
rect 204640 69520 204650 69590
rect 204850 69520 204860 69590
rect 204640 69480 204860 69520
rect 204640 69410 204650 69480
rect 204850 69410 204860 69480
rect 204640 69360 204860 69410
rect 205140 69590 205360 69640
rect 205140 69520 205150 69590
rect 205350 69520 205360 69590
rect 205140 69480 205360 69520
rect 205140 69410 205150 69480
rect 205350 69410 205360 69480
rect 205140 69360 205360 69410
rect 205640 69590 205860 69640
rect 205640 69520 205650 69590
rect 205850 69520 205860 69590
rect 205640 69480 205860 69520
rect 205640 69410 205650 69480
rect 205850 69410 205860 69480
rect 205640 69360 205860 69410
rect 206140 69590 206360 69640
rect 206140 69520 206150 69590
rect 206350 69520 206360 69590
rect 206140 69480 206360 69520
rect 206140 69410 206150 69480
rect 206350 69410 206360 69480
rect 206140 69360 206360 69410
rect 206640 69590 206860 69640
rect 206640 69520 206650 69590
rect 206850 69520 206860 69590
rect 206640 69480 206860 69520
rect 206640 69410 206650 69480
rect 206850 69410 206860 69480
rect 206640 69360 206860 69410
rect 207140 69590 207360 69640
rect 207140 69520 207150 69590
rect 207350 69520 207360 69590
rect 207140 69480 207360 69520
rect 207140 69410 207150 69480
rect 207350 69410 207360 69480
rect 207140 69360 207360 69410
rect 207640 69590 207860 69640
rect 207640 69520 207650 69590
rect 207850 69520 207860 69590
rect 207640 69480 207860 69520
rect 207640 69410 207650 69480
rect 207850 69410 207860 69480
rect 207640 69360 207860 69410
rect 196000 69350 208000 69360
rect 196000 69150 196020 69350
rect 196090 69150 196410 69350
rect 196480 69150 196520 69350
rect 196590 69150 196910 69350
rect 196980 69150 197020 69350
rect 197090 69150 197410 69350
rect 197480 69150 197520 69350
rect 197590 69150 197910 69350
rect 197980 69150 198020 69350
rect 198090 69150 198410 69350
rect 198480 69150 198520 69350
rect 198590 69150 198910 69350
rect 198980 69150 199020 69350
rect 199090 69150 199410 69350
rect 199480 69150 199520 69350
rect 199590 69150 199910 69350
rect 199980 69150 200020 69350
rect 200090 69150 200410 69350
rect 200480 69150 200520 69350
rect 200590 69150 200910 69350
rect 200980 69150 201020 69350
rect 201090 69150 201410 69350
rect 201480 69150 201520 69350
rect 201590 69150 201910 69350
rect 201980 69150 202020 69350
rect 202090 69150 202410 69350
rect 202480 69150 202520 69350
rect 202590 69150 202910 69350
rect 202980 69150 203020 69350
rect 203090 69150 203410 69350
rect 203480 69150 203520 69350
rect 203590 69150 203910 69350
rect 203980 69150 204020 69350
rect 204090 69150 204410 69350
rect 204480 69150 204520 69350
rect 204590 69150 204910 69350
rect 204980 69150 205020 69350
rect 205090 69150 205410 69350
rect 205480 69150 205520 69350
rect 205590 69150 205910 69350
rect 205980 69150 206020 69350
rect 206090 69150 206410 69350
rect 206480 69150 206520 69350
rect 206590 69150 206910 69350
rect 206980 69150 207020 69350
rect 207090 69150 207410 69350
rect 207480 69150 207520 69350
rect 207590 69150 207910 69350
rect 207980 69150 208000 69350
rect 196000 69140 208000 69150
rect 196140 69090 196360 69140
rect 196140 69020 196150 69090
rect 196350 69020 196360 69090
rect 196140 68980 196360 69020
rect 196140 68910 196150 68980
rect 196350 68910 196360 68980
rect 196140 68860 196360 68910
rect 196640 69090 196860 69140
rect 196640 69020 196650 69090
rect 196850 69020 196860 69090
rect 196640 68980 196860 69020
rect 196640 68910 196650 68980
rect 196850 68910 196860 68980
rect 196640 68860 196860 68910
rect 197140 69090 197360 69140
rect 197140 69020 197150 69090
rect 197350 69020 197360 69090
rect 197140 68980 197360 69020
rect 197140 68910 197150 68980
rect 197350 68910 197360 68980
rect 197140 68860 197360 68910
rect 197640 69090 197860 69140
rect 197640 69020 197650 69090
rect 197850 69020 197860 69090
rect 197640 68980 197860 69020
rect 197640 68910 197650 68980
rect 197850 68910 197860 68980
rect 197640 68860 197860 68910
rect 198140 69090 198360 69140
rect 198140 69020 198150 69090
rect 198350 69020 198360 69090
rect 198140 68980 198360 69020
rect 198140 68910 198150 68980
rect 198350 68910 198360 68980
rect 198140 68860 198360 68910
rect 198640 69090 198860 69140
rect 198640 69020 198650 69090
rect 198850 69020 198860 69090
rect 198640 68980 198860 69020
rect 198640 68910 198650 68980
rect 198850 68910 198860 68980
rect 198640 68860 198860 68910
rect 199140 69090 199360 69140
rect 199140 69020 199150 69090
rect 199350 69020 199360 69090
rect 199140 68980 199360 69020
rect 199140 68910 199150 68980
rect 199350 68910 199360 68980
rect 199140 68860 199360 68910
rect 199640 69090 199860 69140
rect 199640 69020 199650 69090
rect 199850 69020 199860 69090
rect 199640 68980 199860 69020
rect 199640 68910 199650 68980
rect 199850 68910 199860 68980
rect 199640 68860 199860 68910
rect 200140 69090 200360 69140
rect 200140 69020 200150 69090
rect 200350 69020 200360 69090
rect 200140 68980 200360 69020
rect 200140 68910 200150 68980
rect 200350 68910 200360 68980
rect 200140 68860 200360 68910
rect 200640 69090 200860 69140
rect 200640 69020 200650 69090
rect 200850 69020 200860 69090
rect 200640 68980 200860 69020
rect 200640 68910 200650 68980
rect 200850 68910 200860 68980
rect 200640 68860 200860 68910
rect 201140 69090 201360 69140
rect 201140 69020 201150 69090
rect 201350 69020 201360 69090
rect 201140 68980 201360 69020
rect 201140 68910 201150 68980
rect 201350 68910 201360 68980
rect 201140 68860 201360 68910
rect 201640 69090 201860 69140
rect 201640 69020 201650 69090
rect 201850 69020 201860 69090
rect 201640 68980 201860 69020
rect 201640 68910 201650 68980
rect 201850 68910 201860 68980
rect 201640 68860 201860 68910
rect 202140 69090 202360 69140
rect 202140 69020 202150 69090
rect 202350 69020 202360 69090
rect 202140 68980 202360 69020
rect 202140 68910 202150 68980
rect 202350 68910 202360 68980
rect 202140 68860 202360 68910
rect 202640 69090 202860 69140
rect 202640 69020 202650 69090
rect 202850 69020 202860 69090
rect 202640 68980 202860 69020
rect 202640 68910 202650 68980
rect 202850 68910 202860 68980
rect 202640 68860 202860 68910
rect 203140 69090 203360 69140
rect 203140 69020 203150 69090
rect 203350 69020 203360 69090
rect 203140 68980 203360 69020
rect 203140 68910 203150 68980
rect 203350 68910 203360 68980
rect 203140 68860 203360 68910
rect 203640 69090 203860 69140
rect 203640 69020 203650 69090
rect 203850 69020 203860 69090
rect 203640 68980 203860 69020
rect 203640 68910 203650 68980
rect 203850 68910 203860 68980
rect 203640 68860 203860 68910
rect 204140 69090 204360 69140
rect 204140 69020 204150 69090
rect 204350 69020 204360 69090
rect 204140 68980 204360 69020
rect 204140 68910 204150 68980
rect 204350 68910 204360 68980
rect 204140 68860 204360 68910
rect 204640 69090 204860 69140
rect 204640 69020 204650 69090
rect 204850 69020 204860 69090
rect 204640 68980 204860 69020
rect 204640 68910 204650 68980
rect 204850 68910 204860 68980
rect 204640 68860 204860 68910
rect 205140 69090 205360 69140
rect 205140 69020 205150 69090
rect 205350 69020 205360 69090
rect 205140 68980 205360 69020
rect 205140 68910 205150 68980
rect 205350 68910 205360 68980
rect 205140 68860 205360 68910
rect 205640 69090 205860 69140
rect 205640 69020 205650 69090
rect 205850 69020 205860 69090
rect 205640 68980 205860 69020
rect 205640 68910 205650 68980
rect 205850 68910 205860 68980
rect 205640 68860 205860 68910
rect 206140 69090 206360 69140
rect 206140 69020 206150 69090
rect 206350 69020 206360 69090
rect 206140 68980 206360 69020
rect 206140 68910 206150 68980
rect 206350 68910 206360 68980
rect 206140 68860 206360 68910
rect 206640 69090 206860 69140
rect 206640 69020 206650 69090
rect 206850 69020 206860 69090
rect 206640 68980 206860 69020
rect 206640 68910 206650 68980
rect 206850 68910 206860 68980
rect 206640 68860 206860 68910
rect 207140 69090 207360 69140
rect 207140 69020 207150 69090
rect 207350 69020 207360 69090
rect 207140 68980 207360 69020
rect 207140 68910 207150 68980
rect 207350 68910 207360 68980
rect 207140 68860 207360 68910
rect 207640 69090 207860 69140
rect 207640 69020 207650 69090
rect 207850 69020 207860 69090
rect 207640 68980 207860 69020
rect 207640 68910 207650 68980
rect 207850 68910 207860 68980
rect 207640 68860 207860 68910
rect 196000 68850 208000 68860
rect 196000 68650 196020 68850
rect 196090 68650 196410 68850
rect 196480 68650 196520 68850
rect 196590 68650 196910 68850
rect 196980 68650 197020 68850
rect 197090 68650 197410 68850
rect 197480 68650 197520 68850
rect 197590 68650 197910 68850
rect 197980 68650 198020 68850
rect 198090 68650 198410 68850
rect 198480 68650 198520 68850
rect 198590 68650 198910 68850
rect 198980 68650 199020 68850
rect 199090 68650 199410 68850
rect 199480 68650 199520 68850
rect 199590 68650 199910 68850
rect 199980 68650 200020 68850
rect 200090 68650 200410 68850
rect 200480 68650 200520 68850
rect 200590 68650 200910 68850
rect 200980 68650 201020 68850
rect 201090 68650 201410 68850
rect 201480 68650 201520 68850
rect 201590 68650 201910 68850
rect 201980 68650 202020 68850
rect 202090 68650 202410 68850
rect 202480 68650 202520 68850
rect 202590 68650 202910 68850
rect 202980 68650 203020 68850
rect 203090 68650 203410 68850
rect 203480 68650 203520 68850
rect 203590 68650 203910 68850
rect 203980 68650 204020 68850
rect 204090 68650 204410 68850
rect 204480 68650 204520 68850
rect 204590 68650 204910 68850
rect 204980 68650 205020 68850
rect 205090 68650 205410 68850
rect 205480 68650 205520 68850
rect 205590 68650 205910 68850
rect 205980 68650 206020 68850
rect 206090 68650 206410 68850
rect 206480 68650 206520 68850
rect 206590 68650 206910 68850
rect 206980 68650 207020 68850
rect 207090 68650 207410 68850
rect 207480 68650 207520 68850
rect 207590 68650 207910 68850
rect 207980 68650 208000 68850
rect 196000 68640 208000 68650
rect 196140 68590 196360 68640
rect 196140 68520 196150 68590
rect 196350 68520 196360 68590
rect 196140 68480 196360 68520
rect 196140 68410 196150 68480
rect 196350 68410 196360 68480
rect 196140 68360 196360 68410
rect 196640 68590 196860 68640
rect 196640 68520 196650 68590
rect 196850 68520 196860 68590
rect 196640 68480 196860 68520
rect 196640 68410 196650 68480
rect 196850 68410 196860 68480
rect 196640 68360 196860 68410
rect 197140 68590 197360 68640
rect 197140 68520 197150 68590
rect 197350 68520 197360 68590
rect 197140 68480 197360 68520
rect 197140 68410 197150 68480
rect 197350 68410 197360 68480
rect 197140 68360 197360 68410
rect 197640 68590 197860 68640
rect 197640 68520 197650 68590
rect 197850 68520 197860 68590
rect 197640 68480 197860 68520
rect 197640 68410 197650 68480
rect 197850 68410 197860 68480
rect 197640 68360 197860 68410
rect 198140 68590 198360 68640
rect 198140 68520 198150 68590
rect 198350 68520 198360 68590
rect 198140 68480 198360 68520
rect 198140 68410 198150 68480
rect 198350 68410 198360 68480
rect 198140 68360 198360 68410
rect 198640 68590 198860 68640
rect 198640 68520 198650 68590
rect 198850 68520 198860 68590
rect 198640 68480 198860 68520
rect 198640 68410 198650 68480
rect 198850 68410 198860 68480
rect 198640 68360 198860 68410
rect 199140 68590 199360 68640
rect 199140 68520 199150 68590
rect 199350 68520 199360 68590
rect 199140 68480 199360 68520
rect 199140 68410 199150 68480
rect 199350 68410 199360 68480
rect 199140 68360 199360 68410
rect 199640 68590 199860 68640
rect 199640 68520 199650 68590
rect 199850 68520 199860 68590
rect 199640 68480 199860 68520
rect 199640 68410 199650 68480
rect 199850 68410 199860 68480
rect 199640 68360 199860 68410
rect 200140 68590 200360 68640
rect 200140 68520 200150 68590
rect 200350 68520 200360 68590
rect 200140 68480 200360 68520
rect 200140 68410 200150 68480
rect 200350 68410 200360 68480
rect 200140 68360 200360 68410
rect 200640 68590 200860 68640
rect 200640 68520 200650 68590
rect 200850 68520 200860 68590
rect 200640 68480 200860 68520
rect 200640 68410 200650 68480
rect 200850 68410 200860 68480
rect 200640 68360 200860 68410
rect 201140 68590 201360 68640
rect 201140 68520 201150 68590
rect 201350 68520 201360 68590
rect 201140 68480 201360 68520
rect 201140 68410 201150 68480
rect 201350 68410 201360 68480
rect 201140 68360 201360 68410
rect 201640 68590 201860 68640
rect 201640 68520 201650 68590
rect 201850 68520 201860 68590
rect 201640 68480 201860 68520
rect 201640 68410 201650 68480
rect 201850 68410 201860 68480
rect 201640 68360 201860 68410
rect 202140 68590 202360 68640
rect 202140 68520 202150 68590
rect 202350 68520 202360 68590
rect 202140 68480 202360 68520
rect 202140 68410 202150 68480
rect 202350 68410 202360 68480
rect 202140 68360 202360 68410
rect 202640 68590 202860 68640
rect 202640 68520 202650 68590
rect 202850 68520 202860 68590
rect 202640 68480 202860 68520
rect 202640 68410 202650 68480
rect 202850 68410 202860 68480
rect 202640 68360 202860 68410
rect 203140 68590 203360 68640
rect 203140 68520 203150 68590
rect 203350 68520 203360 68590
rect 203140 68480 203360 68520
rect 203140 68410 203150 68480
rect 203350 68410 203360 68480
rect 203140 68360 203360 68410
rect 203640 68590 203860 68640
rect 203640 68520 203650 68590
rect 203850 68520 203860 68590
rect 203640 68480 203860 68520
rect 203640 68410 203650 68480
rect 203850 68410 203860 68480
rect 203640 68360 203860 68410
rect 204140 68590 204360 68640
rect 204140 68520 204150 68590
rect 204350 68520 204360 68590
rect 204140 68480 204360 68520
rect 204140 68410 204150 68480
rect 204350 68410 204360 68480
rect 204140 68360 204360 68410
rect 204640 68590 204860 68640
rect 204640 68520 204650 68590
rect 204850 68520 204860 68590
rect 204640 68480 204860 68520
rect 204640 68410 204650 68480
rect 204850 68410 204860 68480
rect 204640 68360 204860 68410
rect 205140 68590 205360 68640
rect 205140 68520 205150 68590
rect 205350 68520 205360 68590
rect 205140 68480 205360 68520
rect 205140 68410 205150 68480
rect 205350 68410 205360 68480
rect 205140 68360 205360 68410
rect 205640 68590 205860 68640
rect 205640 68520 205650 68590
rect 205850 68520 205860 68590
rect 205640 68480 205860 68520
rect 205640 68410 205650 68480
rect 205850 68410 205860 68480
rect 205640 68360 205860 68410
rect 206140 68590 206360 68640
rect 206140 68520 206150 68590
rect 206350 68520 206360 68590
rect 206140 68480 206360 68520
rect 206140 68410 206150 68480
rect 206350 68410 206360 68480
rect 206140 68360 206360 68410
rect 206640 68590 206860 68640
rect 206640 68520 206650 68590
rect 206850 68520 206860 68590
rect 206640 68480 206860 68520
rect 206640 68410 206650 68480
rect 206850 68410 206860 68480
rect 206640 68360 206860 68410
rect 207140 68590 207360 68640
rect 207140 68520 207150 68590
rect 207350 68520 207360 68590
rect 207140 68480 207360 68520
rect 207140 68410 207150 68480
rect 207350 68410 207360 68480
rect 207140 68360 207360 68410
rect 207640 68590 207860 68640
rect 207640 68520 207650 68590
rect 207850 68520 207860 68590
rect 207640 68480 207860 68520
rect 207640 68410 207650 68480
rect 207850 68410 207860 68480
rect 207640 68360 207860 68410
rect 196000 68350 208000 68360
rect 196000 68150 196020 68350
rect 196090 68150 196410 68350
rect 196480 68150 196520 68350
rect 196590 68150 196910 68350
rect 196980 68150 197020 68350
rect 197090 68150 197410 68350
rect 197480 68150 197520 68350
rect 197590 68150 197910 68350
rect 197980 68150 198020 68350
rect 198090 68150 198410 68350
rect 198480 68150 198520 68350
rect 198590 68150 198910 68350
rect 198980 68150 199020 68350
rect 199090 68150 199410 68350
rect 199480 68150 199520 68350
rect 199590 68150 199910 68350
rect 199980 68150 200020 68350
rect 200090 68150 200410 68350
rect 200480 68150 200520 68350
rect 200590 68150 200910 68350
rect 200980 68150 201020 68350
rect 201090 68150 201410 68350
rect 201480 68150 201520 68350
rect 201590 68150 201910 68350
rect 201980 68150 202020 68350
rect 202090 68150 202410 68350
rect 202480 68150 202520 68350
rect 202590 68150 202910 68350
rect 202980 68150 203020 68350
rect 203090 68150 203410 68350
rect 203480 68150 203520 68350
rect 203590 68150 203910 68350
rect 203980 68150 204020 68350
rect 204090 68150 204410 68350
rect 204480 68150 204520 68350
rect 204590 68150 204910 68350
rect 204980 68150 205020 68350
rect 205090 68150 205410 68350
rect 205480 68150 205520 68350
rect 205590 68150 205910 68350
rect 205980 68150 206020 68350
rect 206090 68150 206410 68350
rect 206480 68150 206520 68350
rect 206590 68150 206910 68350
rect 206980 68150 207020 68350
rect 207090 68150 207410 68350
rect 207480 68150 207520 68350
rect 207590 68150 207910 68350
rect 207980 68150 208000 68350
rect 196000 68140 208000 68150
rect 196140 68090 196360 68140
rect 196140 68020 196150 68090
rect 196350 68020 196360 68090
rect 196140 67980 196360 68020
rect 196140 67910 196150 67980
rect 196350 67910 196360 67980
rect 196140 67860 196360 67910
rect 196640 68090 196860 68140
rect 196640 68020 196650 68090
rect 196850 68020 196860 68090
rect 196640 67980 196860 68020
rect 196640 67910 196650 67980
rect 196850 67910 196860 67980
rect 196640 67860 196860 67910
rect 197140 68090 197360 68140
rect 197140 68020 197150 68090
rect 197350 68020 197360 68090
rect 197140 67980 197360 68020
rect 197140 67910 197150 67980
rect 197350 67910 197360 67980
rect 197140 67860 197360 67910
rect 197640 68090 197860 68140
rect 197640 68020 197650 68090
rect 197850 68020 197860 68090
rect 197640 67980 197860 68020
rect 197640 67910 197650 67980
rect 197850 67910 197860 67980
rect 197640 67860 197860 67910
rect 198140 68090 198360 68140
rect 198140 68020 198150 68090
rect 198350 68020 198360 68090
rect 198140 67980 198360 68020
rect 198140 67910 198150 67980
rect 198350 67910 198360 67980
rect 198140 67860 198360 67910
rect 198640 68090 198860 68140
rect 198640 68020 198650 68090
rect 198850 68020 198860 68090
rect 198640 67980 198860 68020
rect 198640 67910 198650 67980
rect 198850 67910 198860 67980
rect 198640 67860 198860 67910
rect 199140 68090 199360 68140
rect 199140 68020 199150 68090
rect 199350 68020 199360 68090
rect 199140 67980 199360 68020
rect 199140 67910 199150 67980
rect 199350 67910 199360 67980
rect 199140 67860 199360 67910
rect 199640 68090 199860 68140
rect 199640 68020 199650 68090
rect 199850 68020 199860 68090
rect 199640 67980 199860 68020
rect 199640 67910 199650 67980
rect 199850 67910 199860 67980
rect 199640 67860 199860 67910
rect 200140 68090 200360 68140
rect 200140 68020 200150 68090
rect 200350 68020 200360 68090
rect 200140 67980 200360 68020
rect 200140 67910 200150 67980
rect 200350 67910 200360 67980
rect 200140 67860 200360 67910
rect 200640 68090 200860 68140
rect 200640 68020 200650 68090
rect 200850 68020 200860 68090
rect 200640 67980 200860 68020
rect 200640 67910 200650 67980
rect 200850 67910 200860 67980
rect 200640 67860 200860 67910
rect 201140 68090 201360 68140
rect 201140 68020 201150 68090
rect 201350 68020 201360 68090
rect 201140 67980 201360 68020
rect 201140 67910 201150 67980
rect 201350 67910 201360 67980
rect 201140 67860 201360 67910
rect 201640 68090 201860 68140
rect 201640 68020 201650 68090
rect 201850 68020 201860 68090
rect 201640 67980 201860 68020
rect 201640 67910 201650 67980
rect 201850 67910 201860 67980
rect 201640 67860 201860 67910
rect 202140 68090 202360 68140
rect 202140 68020 202150 68090
rect 202350 68020 202360 68090
rect 202140 67980 202360 68020
rect 202140 67910 202150 67980
rect 202350 67910 202360 67980
rect 202140 67860 202360 67910
rect 202640 68090 202860 68140
rect 202640 68020 202650 68090
rect 202850 68020 202860 68090
rect 202640 67980 202860 68020
rect 202640 67910 202650 67980
rect 202850 67910 202860 67980
rect 202640 67860 202860 67910
rect 203140 68090 203360 68140
rect 203140 68020 203150 68090
rect 203350 68020 203360 68090
rect 203140 67980 203360 68020
rect 203140 67910 203150 67980
rect 203350 67910 203360 67980
rect 203140 67860 203360 67910
rect 203640 68090 203860 68140
rect 203640 68020 203650 68090
rect 203850 68020 203860 68090
rect 203640 67980 203860 68020
rect 203640 67910 203650 67980
rect 203850 67910 203860 67980
rect 203640 67860 203860 67910
rect 204140 68090 204360 68140
rect 204140 68020 204150 68090
rect 204350 68020 204360 68090
rect 204140 67980 204360 68020
rect 204140 67910 204150 67980
rect 204350 67910 204360 67980
rect 204140 67860 204360 67910
rect 204640 68090 204860 68140
rect 204640 68020 204650 68090
rect 204850 68020 204860 68090
rect 204640 67980 204860 68020
rect 204640 67910 204650 67980
rect 204850 67910 204860 67980
rect 204640 67860 204860 67910
rect 205140 68090 205360 68140
rect 205140 68020 205150 68090
rect 205350 68020 205360 68090
rect 205140 67980 205360 68020
rect 205140 67910 205150 67980
rect 205350 67910 205360 67980
rect 205140 67860 205360 67910
rect 205640 68090 205860 68140
rect 205640 68020 205650 68090
rect 205850 68020 205860 68090
rect 205640 67980 205860 68020
rect 205640 67910 205650 67980
rect 205850 67910 205860 67980
rect 205640 67860 205860 67910
rect 206140 68090 206360 68140
rect 206140 68020 206150 68090
rect 206350 68020 206360 68090
rect 206140 67980 206360 68020
rect 206140 67910 206150 67980
rect 206350 67910 206360 67980
rect 206140 67860 206360 67910
rect 206640 68090 206860 68140
rect 206640 68020 206650 68090
rect 206850 68020 206860 68090
rect 206640 67980 206860 68020
rect 206640 67910 206650 67980
rect 206850 67910 206860 67980
rect 206640 67860 206860 67910
rect 207140 68090 207360 68140
rect 207140 68020 207150 68090
rect 207350 68020 207360 68090
rect 207140 67980 207360 68020
rect 207140 67910 207150 67980
rect 207350 67910 207360 67980
rect 207140 67860 207360 67910
rect 207640 68090 207860 68140
rect 207640 68020 207650 68090
rect 207850 68020 207860 68090
rect 207640 67980 207860 68020
rect 207640 67910 207650 67980
rect 207850 67910 207860 67980
rect 207640 67860 207860 67910
rect 196000 67850 208000 67860
rect 196000 67650 196020 67850
rect 196090 67650 196410 67850
rect 196480 67650 196520 67850
rect 196590 67650 196910 67850
rect 196980 67650 197020 67850
rect 197090 67650 197410 67850
rect 197480 67650 197520 67850
rect 197590 67650 197910 67850
rect 197980 67650 198020 67850
rect 198090 67650 198410 67850
rect 198480 67650 198520 67850
rect 198590 67650 198910 67850
rect 198980 67650 199020 67850
rect 199090 67650 199410 67850
rect 199480 67650 199520 67850
rect 199590 67650 199910 67850
rect 199980 67650 200020 67850
rect 200090 67650 200410 67850
rect 200480 67650 200520 67850
rect 200590 67650 200910 67850
rect 200980 67650 201020 67850
rect 201090 67650 201410 67850
rect 201480 67650 201520 67850
rect 201590 67650 201910 67850
rect 201980 67650 202020 67850
rect 202090 67650 202410 67850
rect 202480 67650 202520 67850
rect 202590 67650 202910 67850
rect 202980 67650 203020 67850
rect 203090 67650 203410 67850
rect 203480 67650 203520 67850
rect 203590 67650 203910 67850
rect 203980 67650 204020 67850
rect 204090 67650 204410 67850
rect 204480 67650 204520 67850
rect 204590 67650 204910 67850
rect 204980 67650 205020 67850
rect 205090 67650 205410 67850
rect 205480 67650 205520 67850
rect 205590 67650 205910 67850
rect 205980 67650 206020 67850
rect 206090 67650 206410 67850
rect 206480 67650 206520 67850
rect 206590 67650 206910 67850
rect 206980 67650 207020 67850
rect 207090 67650 207410 67850
rect 207480 67650 207520 67850
rect 207590 67650 207910 67850
rect 207980 67650 208000 67850
rect 196000 67640 208000 67650
rect 196140 67590 196360 67640
rect 196140 67520 196150 67590
rect 196350 67520 196360 67590
rect 196140 67480 196360 67520
rect 196140 67410 196150 67480
rect 196350 67410 196360 67480
rect 129460 67390 129730 67400
rect 129460 67060 129470 67390
rect 129720 67060 129730 67390
rect 196140 67360 196360 67410
rect 196640 67590 196860 67640
rect 196640 67520 196650 67590
rect 196850 67520 196860 67590
rect 196640 67480 196860 67520
rect 196640 67410 196650 67480
rect 196850 67410 196860 67480
rect 196640 67360 196860 67410
rect 197140 67590 197360 67640
rect 197140 67520 197150 67590
rect 197350 67520 197360 67590
rect 197140 67480 197360 67520
rect 197140 67410 197150 67480
rect 197350 67410 197360 67480
rect 197140 67360 197360 67410
rect 197640 67590 197860 67640
rect 197640 67520 197650 67590
rect 197850 67520 197860 67590
rect 197640 67480 197860 67520
rect 197640 67410 197650 67480
rect 197850 67410 197860 67480
rect 197640 67360 197860 67410
rect 198140 67590 198360 67640
rect 198140 67520 198150 67590
rect 198350 67520 198360 67590
rect 198140 67480 198360 67520
rect 198140 67410 198150 67480
rect 198350 67410 198360 67480
rect 198140 67360 198360 67410
rect 198640 67590 198860 67640
rect 198640 67520 198650 67590
rect 198850 67520 198860 67590
rect 198640 67480 198860 67520
rect 198640 67410 198650 67480
rect 198850 67410 198860 67480
rect 198640 67360 198860 67410
rect 199140 67590 199360 67640
rect 199140 67520 199150 67590
rect 199350 67520 199360 67590
rect 199140 67480 199360 67520
rect 199140 67410 199150 67480
rect 199350 67410 199360 67480
rect 199140 67360 199360 67410
rect 199640 67590 199860 67640
rect 199640 67520 199650 67590
rect 199850 67520 199860 67590
rect 199640 67480 199860 67520
rect 199640 67410 199650 67480
rect 199850 67410 199860 67480
rect 199640 67360 199860 67410
rect 200140 67590 200360 67640
rect 200140 67520 200150 67590
rect 200350 67520 200360 67590
rect 200140 67480 200360 67520
rect 200140 67410 200150 67480
rect 200350 67410 200360 67480
rect 200140 67360 200360 67410
rect 200640 67590 200860 67640
rect 200640 67520 200650 67590
rect 200850 67520 200860 67590
rect 200640 67480 200860 67520
rect 200640 67410 200650 67480
rect 200850 67410 200860 67480
rect 200640 67360 200860 67410
rect 201140 67590 201360 67640
rect 201140 67520 201150 67590
rect 201350 67520 201360 67590
rect 201140 67480 201360 67520
rect 201140 67410 201150 67480
rect 201350 67410 201360 67480
rect 201140 67360 201360 67410
rect 201640 67590 201860 67640
rect 201640 67520 201650 67590
rect 201850 67520 201860 67590
rect 201640 67480 201860 67520
rect 201640 67410 201650 67480
rect 201850 67410 201860 67480
rect 201640 67360 201860 67410
rect 202140 67590 202360 67640
rect 202140 67520 202150 67590
rect 202350 67520 202360 67590
rect 202140 67480 202360 67520
rect 202140 67410 202150 67480
rect 202350 67410 202360 67480
rect 202140 67360 202360 67410
rect 202640 67590 202860 67640
rect 202640 67520 202650 67590
rect 202850 67520 202860 67590
rect 202640 67480 202860 67520
rect 202640 67410 202650 67480
rect 202850 67410 202860 67480
rect 202640 67360 202860 67410
rect 203140 67590 203360 67640
rect 203140 67520 203150 67590
rect 203350 67520 203360 67590
rect 203140 67480 203360 67520
rect 203140 67410 203150 67480
rect 203350 67410 203360 67480
rect 203140 67360 203360 67410
rect 203640 67590 203860 67640
rect 203640 67520 203650 67590
rect 203850 67520 203860 67590
rect 203640 67480 203860 67520
rect 203640 67410 203650 67480
rect 203850 67410 203860 67480
rect 203640 67360 203860 67410
rect 204140 67590 204360 67640
rect 204140 67520 204150 67590
rect 204350 67520 204360 67590
rect 204140 67480 204360 67520
rect 204140 67410 204150 67480
rect 204350 67410 204360 67480
rect 204140 67360 204360 67410
rect 204640 67590 204860 67640
rect 204640 67520 204650 67590
rect 204850 67520 204860 67590
rect 204640 67480 204860 67520
rect 204640 67410 204650 67480
rect 204850 67410 204860 67480
rect 204640 67360 204860 67410
rect 205140 67590 205360 67640
rect 205140 67520 205150 67590
rect 205350 67520 205360 67590
rect 205140 67480 205360 67520
rect 205140 67410 205150 67480
rect 205350 67410 205360 67480
rect 205140 67360 205360 67410
rect 205640 67590 205860 67640
rect 205640 67520 205650 67590
rect 205850 67520 205860 67590
rect 205640 67480 205860 67520
rect 205640 67410 205650 67480
rect 205850 67410 205860 67480
rect 205640 67360 205860 67410
rect 206140 67590 206360 67640
rect 206140 67520 206150 67590
rect 206350 67520 206360 67590
rect 206140 67480 206360 67520
rect 206140 67410 206150 67480
rect 206350 67410 206360 67480
rect 206140 67360 206360 67410
rect 206640 67590 206860 67640
rect 206640 67520 206650 67590
rect 206850 67520 206860 67590
rect 206640 67480 206860 67520
rect 206640 67410 206650 67480
rect 206850 67410 206860 67480
rect 206640 67360 206860 67410
rect 207140 67590 207360 67640
rect 207140 67520 207150 67590
rect 207350 67520 207360 67590
rect 207140 67480 207360 67520
rect 207140 67410 207150 67480
rect 207350 67410 207360 67480
rect 207140 67360 207360 67410
rect 207640 67590 207860 67640
rect 207640 67520 207650 67590
rect 207850 67520 207860 67590
rect 207640 67480 207860 67520
rect 207640 67410 207650 67480
rect 207850 67410 207860 67480
rect 207640 67360 207860 67410
rect 196000 67350 208000 67360
rect 196000 67150 196020 67350
rect 196090 67150 196410 67350
rect 196480 67150 196520 67350
rect 196590 67150 196910 67350
rect 196980 67150 197020 67350
rect 197090 67150 197410 67350
rect 197480 67150 197520 67350
rect 197590 67150 197910 67350
rect 197980 67150 198020 67350
rect 198090 67150 198410 67350
rect 198480 67150 198520 67350
rect 198590 67150 198910 67350
rect 198980 67150 199020 67350
rect 199090 67150 199410 67350
rect 199480 67150 199520 67350
rect 199590 67150 199910 67350
rect 199980 67150 200020 67350
rect 200090 67150 200410 67350
rect 200480 67150 200520 67350
rect 200590 67150 200910 67350
rect 200980 67150 201020 67350
rect 201090 67150 201410 67350
rect 201480 67150 201520 67350
rect 201590 67150 201910 67350
rect 201980 67150 202020 67350
rect 202090 67150 202410 67350
rect 202480 67150 202520 67350
rect 202590 67150 202910 67350
rect 202980 67150 203020 67350
rect 203090 67150 203410 67350
rect 203480 67150 203520 67350
rect 203590 67150 203910 67350
rect 203980 67150 204020 67350
rect 204090 67150 204410 67350
rect 204480 67150 204520 67350
rect 204590 67150 204910 67350
rect 204980 67150 205020 67350
rect 205090 67150 205410 67350
rect 205480 67150 205520 67350
rect 205590 67150 205910 67350
rect 205980 67150 206020 67350
rect 206090 67150 206410 67350
rect 206480 67150 206520 67350
rect 206590 67150 206910 67350
rect 206980 67150 207020 67350
rect 207090 67150 207410 67350
rect 207480 67150 207520 67350
rect 207590 67150 207910 67350
rect 207980 67150 208000 67350
rect 196000 67140 208000 67150
rect 129460 67050 129730 67060
rect 129590 66950 129730 67050
rect 196140 67090 196360 67140
rect 196140 67020 196150 67090
rect 196350 67020 196360 67090
rect 196140 66980 196360 67020
rect 129590 66850 137560 66950
rect 196140 66910 196150 66980
rect 196350 66910 196360 66980
rect 196140 66860 196360 66910
rect 196640 67090 196860 67140
rect 196640 67020 196650 67090
rect 196850 67020 196860 67090
rect 196640 66980 196860 67020
rect 196640 66910 196650 66980
rect 196850 66910 196860 66980
rect 196640 66860 196860 66910
rect 197140 67090 197360 67140
rect 197140 67020 197150 67090
rect 197350 67020 197360 67090
rect 197140 66980 197360 67020
rect 197140 66910 197150 66980
rect 197350 66910 197360 66980
rect 197140 66860 197360 66910
rect 197640 67090 197860 67140
rect 197640 67020 197650 67090
rect 197850 67020 197860 67090
rect 197640 66980 197860 67020
rect 197640 66910 197650 66980
rect 197850 66910 197860 66980
rect 197640 66860 197860 66910
rect 198140 67090 198360 67140
rect 198140 67020 198150 67090
rect 198350 67020 198360 67090
rect 198140 66980 198360 67020
rect 198140 66910 198150 66980
rect 198350 66910 198360 66980
rect 198140 66860 198360 66910
rect 198640 67090 198860 67140
rect 198640 67020 198650 67090
rect 198850 67020 198860 67090
rect 198640 66980 198860 67020
rect 198640 66910 198650 66980
rect 198850 66910 198860 66980
rect 198640 66860 198860 66910
rect 199140 67090 199360 67140
rect 199140 67020 199150 67090
rect 199350 67020 199360 67090
rect 199140 66980 199360 67020
rect 199140 66910 199150 66980
rect 199350 66910 199360 66980
rect 199140 66860 199360 66910
rect 199640 67090 199860 67140
rect 199640 67020 199650 67090
rect 199850 67020 199860 67090
rect 199640 66980 199860 67020
rect 199640 66910 199650 66980
rect 199850 66910 199860 66980
rect 199640 66860 199860 66910
rect 200140 67090 200360 67140
rect 200140 67020 200150 67090
rect 200350 67020 200360 67090
rect 200140 66980 200360 67020
rect 200140 66910 200150 66980
rect 200350 66910 200360 66980
rect 200140 66860 200360 66910
rect 200640 67090 200860 67140
rect 200640 67020 200650 67090
rect 200850 67020 200860 67090
rect 200640 66980 200860 67020
rect 200640 66910 200650 66980
rect 200850 66910 200860 66980
rect 200640 66860 200860 66910
rect 201140 67090 201360 67140
rect 201140 67020 201150 67090
rect 201350 67020 201360 67090
rect 201140 66980 201360 67020
rect 201140 66910 201150 66980
rect 201350 66910 201360 66980
rect 201140 66860 201360 66910
rect 201640 67090 201860 67140
rect 201640 67020 201650 67090
rect 201850 67020 201860 67090
rect 201640 66980 201860 67020
rect 201640 66910 201650 66980
rect 201850 66910 201860 66980
rect 201640 66860 201860 66910
rect 202140 67090 202360 67140
rect 202140 67020 202150 67090
rect 202350 67020 202360 67090
rect 202140 66980 202360 67020
rect 202140 66910 202150 66980
rect 202350 66910 202360 66980
rect 202140 66860 202360 66910
rect 202640 67090 202860 67140
rect 202640 67020 202650 67090
rect 202850 67020 202860 67090
rect 202640 66980 202860 67020
rect 202640 66910 202650 66980
rect 202850 66910 202860 66980
rect 202640 66860 202860 66910
rect 203140 67090 203360 67140
rect 203140 67020 203150 67090
rect 203350 67020 203360 67090
rect 203140 66980 203360 67020
rect 203140 66910 203150 66980
rect 203350 66910 203360 66980
rect 203140 66860 203360 66910
rect 203640 67090 203860 67140
rect 203640 67020 203650 67090
rect 203850 67020 203860 67090
rect 203640 66980 203860 67020
rect 203640 66910 203650 66980
rect 203850 66910 203860 66980
rect 203640 66860 203860 66910
rect 204140 67090 204360 67140
rect 204140 67020 204150 67090
rect 204350 67020 204360 67090
rect 204140 66980 204360 67020
rect 204140 66910 204150 66980
rect 204350 66910 204360 66980
rect 204140 66860 204360 66910
rect 204640 67090 204860 67140
rect 204640 67020 204650 67090
rect 204850 67020 204860 67090
rect 204640 66980 204860 67020
rect 204640 66910 204650 66980
rect 204850 66910 204860 66980
rect 204640 66860 204860 66910
rect 205140 67090 205360 67140
rect 205140 67020 205150 67090
rect 205350 67020 205360 67090
rect 205140 66980 205360 67020
rect 205140 66910 205150 66980
rect 205350 66910 205360 66980
rect 205140 66860 205360 66910
rect 205640 67090 205860 67140
rect 205640 67020 205650 67090
rect 205850 67020 205860 67090
rect 205640 66980 205860 67020
rect 205640 66910 205650 66980
rect 205850 66910 205860 66980
rect 205640 66860 205860 66910
rect 206140 67090 206360 67140
rect 206140 67020 206150 67090
rect 206350 67020 206360 67090
rect 206140 66980 206360 67020
rect 206140 66910 206150 66980
rect 206350 66910 206360 66980
rect 206140 66860 206360 66910
rect 206640 67090 206860 67140
rect 206640 67020 206650 67090
rect 206850 67020 206860 67090
rect 206640 66980 206860 67020
rect 206640 66910 206650 66980
rect 206850 66910 206860 66980
rect 206640 66860 206860 66910
rect 207140 67090 207360 67140
rect 207140 67020 207150 67090
rect 207350 67020 207360 67090
rect 207140 66980 207360 67020
rect 207140 66910 207150 66980
rect 207350 66910 207360 66980
rect 207140 66860 207360 66910
rect 207640 67090 207860 67140
rect 207640 67020 207650 67090
rect 207850 67020 207860 67090
rect 207640 66980 207860 67020
rect 207640 66910 207650 66980
rect 207850 66910 207860 66980
rect 207640 66860 207860 66910
rect 137460 66110 137560 66850
rect 196000 66850 208000 66860
rect 196000 66650 196020 66850
rect 196090 66650 196410 66850
rect 196480 66650 196520 66850
rect 196590 66650 196910 66850
rect 196980 66650 197020 66850
rect 197090 66650 197410 66850
rect 197480 66650 197520 66850
rect 197590 66650 197910 66850
rect 197980 66650 198020 66850
rect 198090 66650 198410 66850
rect 198480 66650 198520 66850
rect 198590 66650 198910 66850
rect 198980 66650 199020 66850
rect 199090 66650 199410 66850
rect 199480 66650 199520 66850
rect 199590 66650 199910 66850
rect 199980 66650 200020 66850
rect 200090 66650 200410 66850
rect 200480 66650 200520 66850
rect 200590 66650 200910 66850
rect 200980 66650 201020 66850
rect 201090 66650 201410 66850
rect 201480 66650 201520 66850
rect 201590 66650 201910 66850
rect 201980 66650 202020 66850
rect 202090 66650 202410 66850
rect 202480 66650 202520 66850
rect 202590 66650 202910 66850
rect 202980 66650 203020 66850
rect 203090 66650 203410 66850
rect 203480 66650 203520 66850
rect 203590 66650 203910 66850
rect 203980 66650 204020 66850
rect 204090 66650 204410 66850
rect 204480 66650 204520 66850
rect 204590 66650 204910 66850
rect 204980 66650 205020 66850
rect 205090 66650 205410 66850
rect 205480 66650 205520 66850
rect 205590 66650 205910 66850
rect 205980 66650 206020 66850
rect 206090 66650 206410 66850
rect 206480 66650 206520 66850
rect 206590 66650 206910 66850
rect 206980 66650 207020 66850
rect 207090 66650 207410 66850
rect 207480 66650 207520 66850
rect 207590 66650 207910 66850
rect 207980 66650 208000 66850
rect 196000 66640 208000 66650
rect 196140 66590 196360 66640
rect 196140 66520 196150 66590
rect 196350 66520 196360 66590
rect 196140 66480 196360 66520
rect 196140 66410 196150 66480
rect 196350 66410 196360 66480
rect 196140 66360 196360 66410
rect 196640 66590 196860 66640
rect 196640 66520 196650 66590
rect 196850 66520 196860 66590
rect 196640 66480 196860 66520
rect 196640 66410 196650 66480
rect 196850 66410 196860 66480
rect 196640 66360 196860 66410
rect 197140 66590 197360 66640
rect 197140 66520 197150 66590
rect 197350 66520 197360 66590
rect 197140 66480 197360 66520
rect 197140 66410 197150 66480
rect 197350 66410 197360 66480
rect 197140 66360 197360 66410
rect 197640 66590 197860 66640
rect 197640 66520 197650 66590
rect 197850 66520 197860 66590
rect 197640 66480 197860 66520
rect 197640 66410 197650 66480
rect 197850 66410 197860 66480
rect 197640 66360 197860 66410
rect 198140 66590 198360 66640
rect 198140 66520 198150 66590
rect 198350 66520 198360 66590
rect 198140 66480 198360 66520
rect 198140 66410 198150 66480
rect 198350 66410 198360 66480
rect 198140 66360 198360 66410
rect 198640 66590 198860 66640
rect 198640 66520 198650 66590
rect 198850 66520 198860 66590
rect 198640 66480 198860 66520
rect 198640 66410 198650 66480
rect 198850 66410 198860 66480
rect 198640 66360 198860 66410
rect 199140 66590 199360 66640
rect 199140 66520 199150 66590
rect 199350 66520 199360 66590
rect 199140 66480 199360 66520
rect 199140 66410 199150 66480
rect 199350 66410 199360 66480
rect 199140 66360 199360 66410
rect 199640 66590 199860 66640
rect 199640 66520 199650 66590
rect 199850 66520 199860 66590
rect 199640 66480 199860 66520
rect 199640 66410 199650 66480
rect 199850 66410 199860 66480
rect 199640 66360 199860 66410
rect 200140 66590 200360 66640
rect 200140 66520 200150 66590
rect 200350 66520 200360 66590
rect 200140 66480 200360 66520
rect 200140 66410 200150 66480
rect 200350 66410 200360 66480
rect 200140 66360 200360 66410
rect 200640 66590 200860 66640
rect 200640 66520 200650 66590
rect 200850 66520 200860 66590
rect 200640 66480 200860 66520
rect 200640 66410 200650 66480
rect 200850 66410 200860 66480
rect 200640 66360 200860 66410
rect 201140 66590 201360 66640
rect 201140 66520 201150 66590
rect 201350 66520 201360 66590
rect 201140 66480 201360 66520
rect 201140 66410 201150 66480
rect 201350 66410 201360 66480
rect 201140 66360 201360 66410
rect 201640 66590 201860 66640
rect 201640 66520 201650 66590
rect 201850 66520 201860 66590
rect 201640 66480 201860 66520
rect 201640 66410 201650 66480
rect 201850 66410 201860 66480
rect 201640 66360 201860 66410
rect 202140 66590 202360 66640
rect 202140 66520 202150 66590
rect 202350 66520 202360 66590
rect 202140 66480 202360 66520
rect 202140 66410 202150 66480
rect 202350 66410 202360 66480
rect 202140 66360 202360 66410
rect 202640 66590 202860 66640
rect 202640 66520 202650 66590
rect 202850 66520 202860 66590
rect 202640 66480 202860 66520
rect 202640 66410 202650 66480
rect 202850 66410 202860 66480
rect 202640 66360 202860 66410
rect 203140 66590 203360 66640
rect 203140 66520 203150 66590
rect 203350 66520 203360 66590
rect 203140 66480 203360 66520
rect 203140 66410 203150 66480
rect 203350 66410 203360 66480
rect 203140 66360 203360 66410
rect 203640 66590 203860 66640
rect 203640 66520 203650 66590
rect 203850 66520 203860 66590
rect 203640 66480 203860 66520
rect 203640 66410 203650 66480
rect 203850 66410 203860 66480
rect 203640 66360 203860 66410
rect 204140 66590 204360 66640
rect 204140 66520 204150 66590
rect 204350 66520 204360 66590
rect 204140 66480 204360 66520
rect 204140 66410 204150 66480
rect 204350 66410 204360 66480
rect 204140 66360 204360 66410
rect 204640 66590 204860 66640
rect 204640 66520 204650 66590
rect 204850 66520 204860 66590
rect 204640 66480 204860 66520
rect 204640 66410 204650 66480
rect 204850 66410 204860 66480
rect 204640 66360 204860 66410
rect 205140 66590 205360 66640
rect 205140 66520 205150 66590
rect 205350 66520 205360 66590
rect 205140 66480 205360 66520
rect 205140 66410 205150 66480
rect 205350 66410 205360 66480
rect 205140 66360 205360 66410
rect 205640 66590 205860 66640
rect 205640 66520 205650 66590
rect 205850 66520 205860 66590
rect 205640 66480 205860 66520
rect 205640 66410 205650 66480
rect 205850 66410 205860 66480
rect 205640 66360 205860 66410
rect 206140 66590 206360 66640
rect 206140 66520 206150 66590
rect 206350 66520 206360 66590
rect 206140 66480 206360 66520
rect 206140 66410 206150 66480
rect 206350 66410 206360 66480
rect 206140 66360 206360 66410
rect 206640 66590 206860 66640
rect 206640 66520 206650 66590
rect 206850 66520 206860 66590
rect 206640 66480 206860 66520
rect 206640 66410 206650 66480
rect 206850 66410 206860 66480
rect 206640 66360 206860 66410
rect 207140 66590 207360 66640
rect 207140 66520 207150 66590
rect 207350 66520 207360 66590
rect 207140 66480 207360 66520
rect 207140 66410 207150 66480
rect 207350 66410 207360 66480
rect 207140 66360 207360 66410
rect 207640 66590 207860 66640
rect 207640 66520 207650 66590
rect 207850 66520 207860 66590
rect 207640 66480 207860 66520
rect 207640 66410 207650 66480
rect 207850 66410 207860 66480
rect 207640 66360 207860 66410
rect 196000 66350 208000 66360
rect 196000 66150 196020 66350
rect 196090 66150 196410 66350
rect 196480 66150 196520 66350
rect 196590 66150 196910 66350
rect 196980 66150 197020 66350
rect 197090 66150 197410 66350
rect 197480 66150 197520 66350
rect 197590 66150 197910 66350
rect 197980 66150 198020 66350
rect 198090 66150 198410 66350
rect 198480 66150 198520 66350
rect 198590 66150 198910 66350
rect 198980 66150 199020 66350
rect 199090 66150 199410 66350
rect 199480 66150 199520 66350
rect 199590 66150 199910 66350
rect 199980 66150 200020 66350
rect 200090 66150 200410 66350
rect 200480 66150 200520 66350
rect 200590 66150 200910 66350
rect 200980 66150 201020 66350
rect 201090 66150 201410 66350
rect 201480 66150 201520 66350
rect 201590 66150 201910 66350
rect 201980 66150 202020 66350
rect 202090 66150 202410 66350
rect 202480 66150 202520 66350
rect 202590 66150 202910 66350
rect 202980 66150 203020 66350
rect 203090 66150 203410 66350
rect 203480 66150 203520 66350
rect 203590 66150 203910 66350
rect 203980 66150 204020 66350
rect 204090 66150 204410 66350
rect 204480 66150 204520 66350
rect 204590 66150 204910 66350
rect 204980 66150 205020 66350
rect 205090 66150 205410 66350
rect 205480 66150 205520 66350
rect 205590 66150 205910 66350
rect 205980 66150 206020 66350
rect 206090 66150 206410 66350
rect 206480 66150 206520 66350
rect 206590 66150 206910 66350
rect 206980 66150 207020 66350
rect 207090 66150 207410 66350
rect 207480 66150 207520 66350
rect 207590 66150 207910 66350
rect 207980 66150 208000 66350
rect 196000 66140 208000 66150
rect 196140 66090 196360 66140
rect 196140 66020 196150 66090
rect 196350 66020 196360 66090
rect 190140 65980 190360 66000
rect 190140 65910 190150 65980
rect 190350 65910 190360 65980
rect 190140 65860 190360 65910
rect 190640 65980 190860 66000
rect 190640 65910 190650 65980
rect 190850 65910 190860 65980
rect 190640 65860 190860 65910
rect 191140 65980 191360 66000
rect 191140 65910 191150 65980
rect 191350 65910 191360 65980
rect 191140 65860 191360 65910
rect 191640 65980 191860 66000
rect 191640 65910 191650 65980
rect 191850 65910 191860 65980
rect 191640 65860 191860 65910
rect 192140 65980 192360 66000
rect 192140 65910 192150 65980
rect 192350 65910 192360 65980
rect 192140 65860 192360 65910
rect 192640 65980 192860 66000
rect 192640 65910 192650 65980
rect 192850 65910 192860 65980
rect 192640 65860 192860 65910
rect 193140 65980 193360 66000
rect 193140 65910 193150 65980
rect 193350 65910 193360 65980
rect 193140 65860 193360 65910
rect 193640 65980 193860 66000
rect 193640 65910 193650 65980
rect 193850 65910 193860 65980
rect 193640 65860 193860 65910
rect 194140 65980 194360 66000
rect 194140 65910 194150 65980
rect 194350 65910 194360 65980
rect 194140 65860 194360 65910
rect 194640 65980 194860 66000
rect 194640 65910 194650 65980
rect 194850 65910 194860 65980
rect 194640 65860 194860 65910
rect 195140 65980 195360 66000
rect 195140 65910 195150 65980
rect 195350 65910 195360 65980
rect 195140 65860 195360 65910
rect 195640 65980 195860 66000
rect 195640 65910 195650 65980
rect 195850 65910 195860 65980
rect 195640 65860 195860 65910
rect 196140 65980 196360 66020
rect 196140 65910 196150 65980
rect 196350 65910 196360 65980
rect 196140 65860 196360 65910
rect 196640 66090 196860 66140
rect 196640 66020 196650 66090
rect 196850 66020 196860 66090
rect 196640 65980 196860 66020
rect 196640 65910 196650 65980
rect 196850 65910 196860 65980
rect 196640 65860 196860 65910
rect 197140 66090 197360 66140
rect 197140 66020 197150 66090
rect 197350 66020 197360 66090
rect 197140 65980 197360 66020
rect 197140 65910 197150 65980
rect 197350 65910 197360 65980
rect 197140 65860 197360 65910
rect 197640 66090 197860 66140
rect 197640 66020 197650 66090
rect 197850 66020 197860 66090
rect 197640 65980 197860 66020
rect 197640 65910 197650 65980
rect 197850 65910 197860 65980
rect 197640 65860 197860 65910
rect 198140 66090 198360 66140
rect 198140 66020 198150 66090
rect 198350 66020 198360 66090
rect 198140 65980 198360 66020
rect 198140 65910 198150 65980
rect 198350 65910 198360 65980
rect 198140 65860 198360 65910
rect 198640 66090 198860 66140
rect 198640 66020 198650 66090
rect 198850 66020 198860 66090
rect 198640 65980 198860 66020
rect 198640 65910 198650 65980
rect 198850 65910 198860 65980
rect 198640 65860 198860 65910
rect 199140 66090 199360 66140
rect 199140 66020 199150 66090
rect 199350 66020 199360 66090
rect 199140 65980 199360 66020
rect 199140 65910 199150 65980
rect 199350 65910 199360 65980
rect 199140 65860 199360 65910
rect 199640 66090 199860 66140
rect 199640 66020 199650 66090
rect 199850 66020 199860 66090
rect 199640 65980 199860 66020
rect 199640 65910 199650 65980
rect 199850 65910 199860 65980
rect 199640 65860 199860 65910
rect 200140 66090 200360 66140
rect 200140 66020 200150 66090
rect 200350 66020 200360 66090
rect 200140 65980 200360 66020
rect 200140 65910 200150 65980
rect 200350 65910 200360 65980
rect 200140 65860 200360 65910
rect 200640 66090 200860 66140
rect 200640 66020 200650 66090
rect 200850 66020 200860 66090
rect 200640 65980 200860 66020
rect 200640 65910 200650 65980
rect 200850 65910 200860 65980
rect 200640 65860 200860 65910
rect 201140 66090 201360 66140
rect 201140 66020 201150 66090
rect 201350 66020 201360 66090
rect 201140 65980 201360 66020
rect 201140 65910 201150 65980
rect 201350 65910 201360 65980
rect 201140 65860 201360 65910
rect 201640 66090 201860 66140
rect 201640 66020 201650 66090
rect 201850 66020 201860 66090
rect 201640 65980 201860 66020
rect 201640 65910 201650 65980
rect 201850 65910 201860 65980
rect 201640 65860 201860 65910
rect 202140 66090 202360 66140
rect 202140 66020 202150 66090
rect 202350 66020 202360 66090
rect 202140 65980 202360 66020
rect 202140 65910 202150 65980
rect 202350 65910 202360 65980
rect 202140 65860 202360 65910
rect 202640 66090 202860 66140
rect 202640 66020 202650 66090
rect 202850 66020 202860 66090
rect 202640 65980 202860 66020
rect 202640 65910 202650 65980
rect 202850 65910 202860 65980
rect 202640 65860 202860 65910
rect 203140 66090 203360 66140
rect 203140 66020 203150 66090
rect 203350 66020 203360 66090
rect 203140 65980 203360 66020
rect 203140 65910 203150 65980
rect 203350 65910 203360 65980
rect 203140 65860 203360 65910
rect 203640 66090 203860 66140
rect 203640 66020 203650 66090
rect 203850 66020 203860 66090
rect 203640 65980 203860 66020
rect 203640 65910 203650 65980
rect 203850 65910 203860 65980
rect 203640 65860 203860 65910
rect 204140 66090 204360 66140
rect 204140 66020 204150 66090
rect 204350 66020 204360 66090
rect 204140 65980 204360 66020
rect 204140 65910 204150 65980
rect 204350 65910 204360 65980
rect 204140 65860 204360 65910
rect 204640 66090 204860 66140
rect 204640 66020 204650 66090
rect 204850 66020 204860 66090
rect 204640 65980 204860 66020
rect 204640 65910 204650 65980
rect 204850 65910 204860 65980
rect 204640 65860 204860 65910
rect 205140 66090 205360 66140
rect 205140 66020 205150 66090
rect 205350 66020 205360 66090
rect 205140 65980 205360 66020
rect 205140 65910 205150 65980
rect 205350 65910 205360 65980
rect 205140 65860 205360 65910
rect 205640 66090 205860 66140
rect 205640 66020 205650 66090
rect 205850 66020 205860 66090
rect 205640 65980 205860 66020
rect 205640 65910 205650 65980
rect 205850 65910 205860 65980
rect 205640 65860 205860 65910
rect 206140 66090 206360 66140
rect 206140 66020 206150 66090
rect 206350 66020 206360 66090
rect 206140 65980 206360 66020
rect 206140 65910 206150 65980
rect 206350 65910 206360 65980
rect 206140 65860 206360 65910
rect 206640 66090 206860 66140
rect 206640 66020 206650 66090
rect 206850 66020 206860 66090
rect 206640 65980 206860 66020
rect 206640 65910 206650 65980
rect 206850 65910 206860 65980
rect 206640 65860 206860 65910
rect 207140 66090 207360 66140
rect 207140 66020 207150 66090
rect 207350 66020 207360 66090
rect 207140 65980 207360 66020
rect 207140 65910 207150 65980
rect 207350 65910 207360 65980
rect 207140 65860 207360 65910
rect 207640 66090 207860 66140
rect 207640 66020 207650 66090
rect 207850 66020 207860 66090
rect 207640 65980 207860 66020
rect 207640 65910 207650 65980
rect 207850 65910 207860 65980
rect 207640 65860 207860 65910
rect 190000 65850 208000 65860
rect 190000 65650 190020 65850
rect 190090 65650 190410 65850
rect 190480 65650 190520 65850
rect 190590 65650 190910 65850
rect 190980 65650 191020 65850
rect 191090 65650 191410 65850
rect 191480 65650 191520 65850
rect 191590 65650 191910 65850
rect 191980 65650 192020 65850
rect 192090 65650 192410 65850
rect 192480 65650 192520 65850
rect 192590 65650 192910 65850
rect 192980 65650 193020 65850
rect 193090 65650 193410 65850
rect 193480 65650 193520 65850
rect 193590 65650 193910 65850
rect 193980 65650 194020 65850
rect 194090 65650 194410 65850
rect 194480 65650 194520 65850
rect 194590 65650 194910 65850
rect 194980 65650 195020 65850
rect 195090 65650 195410 65850
rect 195480 65650 195520 65850
rect 195590 65650 195910 65850
rect 195980 65650 196020 65850
rect 196090 65650 196410 65850
rect 196480 65650 196520 65850
rect 196590 65650 196910 65850
rect 196980 65650 197020 65850
rect 197090 65650 197410 65850
rect 197480 65650 197520 65850
rect 197590 65650 197910 65850
rect 197980 65650 198020 65850
rect 198090 65650 198410 65850
rect 198480 65650 198520 65850
rect 198590 65650 198910 65850
rect 198980 65650 199020 65850
rect 199090 65650 199410 65850
rect 199480 65650 199520 65850
rect 199590 65650 199910 65850
rect 199980 65650 200020 65850
rect 200090 65650 200410 65850
rect 200480 65650 200520 65850
rect 200590 65650 200910 65850
rect 200980 65650 201020 65850
rect 201090 65650 201410 65850
rect 201480 65650 201520 65850
rect 201590 65650 201910 65850
rect 201980 65650 202020 65850
rect 202090 65650 202410 65850
rect 202480 65650 202520 65850
rect 202590 65650 202910 65850
rect 202980 65650 203020 65850
rect 203090 65650 203410 65850
rect 203480 65650 203520 65850
rect 203590 65650 203910 65850
rect 203980 65650 204020 65850
rect 204090 65650 204410 65850
rect 204480 65650 204520 65850
rect 204590 65650 204910 65850
rect 204980 65650 205020 65850
rect 205090 65650 205410 65850
rect 205480 65650 205520 65850
rect 205590 65650 205910 65850
rect 205980 65650 206020 65850
rect 206090 65650 206410 65850
rect 206480 65650 206520 65850
rect 206590 65650 206910 65850
rect 206980 65650 207020 65850
rect 207090 65650 207410 65850
rect 207480 65650 207520 65850
rect 207590 65650 207910 65850
rect 207980 65650 208000 65850
rect 190000 65640 208000 65650
rect 190140 65590 190360 65640
rect 190140 65520 190150 65590
rect 190350 65520 190360 65590
rect 190140 65480 190360 65520
rect 190140 65410 190150 65480
rect 190350 65410 190360 65480
rect 190140 65360 190360 65410
rect 190640 65590 190860 65640
rect 190640 65520 190650 65590
rect 190850 65520 190860 65590
rect 190640 65480 190860 65520
rect 190640 65410 190650 65480
rect 190850 65410 190860 65480
rect 190640 65360 190860 65410
rect 191140 65590 191360 65640
rect 191140 65520 191150 65590
rect 191350 65520 191360 65590
rect 191140 65480 191360 65520
rect 191140 65410 191150 65480
rect 191350 65410 191360 65480
rect 191140 65360 191360 65410
rect 191640 65590 191860 65640
rect 191640 65520 191650 65590
rect 191850 65520 191860 65590
rect 191640 65480 191860 65520
rect 191640 65410 191650 65480
rect 191850 65410 191860 65480
rect 191640 65360 191860 65410
rect 192140 65590 192360 65640
rect 192140 65520 192150 65590
rect 192350 65520 192360 65590
rect 192140 65480 192360 65520
rect 192140 65410 192150 65480
rect 192350 65410 192360 65480
rect 192140 65360 192360 65410
rect 192640 65590 192860 65640
rect 192640 65520 192650 65590
rect 192850 65520 192860 65590
rect 192640 65480 192860 65520
rect 192640 65410 192650 65480
rect 192850 65410 192860 65480
rect 192640 65360 192860 65410
rect 193140 65590 193360 65640
rect 193140 65520 193150 65590
rect 193350 65520 193360 65590
rect 193140 65480 193360 65520
rect 193140 65410 193150 65480
rect 193350 65410 193360 65480
rect 193140 65360 193360 65410
rect 193640 65590 193860 65640
rect 193640 65520 193650 65590
rect 193850 65520 193860 65590
rect 193640 65480 193860 65520
rect 193640 65410 193650 65480
rect 193850 65410 193860 65480
rect 193640 65360 193860 65410
rect 194140 65590 194360 65640
rect 194140 65520 194150 65590
rect 194350 65520 194360 65590
rect 194140 65480 194360 65520
rect 194140 65410 194150 65480
rect 194350 65410 194360 65480
rect 194140 65360 194360 65410
rect 194640 65590 194860 65640
rect 194640 65520 194650 65590
rect 194850 65520 194860 65590
rect 194640 65480 194860 65520
rect 194640 65410 194650 65480
rect 194850 65410 194860 65480
rect 194640 65360 194860 65410
rect 195140 65590 195360 65640
rect 195140 65520 195150 65590
rect 195350 65520 195360 65590
rect 195140 65480 195360 65520
rect 195140 65410 195150 65480
rect 195350 65410 195360 65480
rect 195140 65360 195360 65410
rect 195640 65590 195860 65640
rect 195640 65520 195650 65590
rect 195850 65520 195860 65590
rect 195640 65480 195860 65520
rect 195640 65410 195650 65480
rect 195850 65410 195860 65480
rect 195640 65360 195860 65410
rect 196140 65590 196360 65640
rect 196140 65520 196150 65590
rect 196350 65520 196360 65590
rect 196140 65480 196360 65520
rect 196140 65410 196150 65480
rect 196350 65410 196360 65480
rect 196140 65360 196360 65410
rect 196640 65590 196860 65640
rect 196640 65520 196650 65590
rect 196850 65520 196860 65590
rect 196640 65480 196860 65520
rect 196640 65410 196650 65480
rect 196850 65410 196860 65480
rect 196640 65360 196860 65410
rect 197140 65590 197360 65640
rect 197140 65520 197150 65590
rect 197350 65520 197360 65590
rect 197140 65480 197360 65520
rect 197140 65410 197150 65480
rect 197350 65410 197360 65480
rect 197140 65360 197360 65410
rect 197640 65590 197860 65640
rect 197640 65520 197650 65590
rect 197850 65520 197860 65590
rect 197640 65480 197860 65520
rect 197640 65410 197650 65480
rect 197850 65410 197860 65480
rect 197640 65360 197860 65410
rect 198140 65590 198360 65640
rect 198140 65520 198150 65590
rect 198350 65520 198360 65590
rect 198140 65480 198360 65520
rect 198140 65410 198150 65480
rect 198350 65410 198360 65480
rect 198140 65360 198360 65410
rect 198640 65590 198860 65640
rect 198640 65520 198650 65590
rect 198850 65520 198860 65590
rect 198640 65480 198860 65520
rect 198640 65410 198650 65480
rect 198850 65410 198860 65480
rect 198640 65360 198860 65410
rect 199140 65590 199360 65640
rect 199140 65520 199150 65590
rect 199350 65520 199360 65590
rect 199140 65480 199360 65520
rect 199140 65410 199150 65480
rect 199350 65410 199360 65480
rect 199140 65360 199360 65410
rect 199640 65590 199860 65640
rect 199640 65520 199650 65590
rect 199850 65520 199860 65590
rect 199640 65480 199860 65520
rect 199640 65410 199650 65480
rect 199850 65410 199860 65480
rect 199640 65360 199860 65410
rect 200140 65590 200360 65640
rect 200140 65520 200150 65590
rect 200350 65520 200360 65590
rect 200140 65480 200360 65520
rect 200140 65410 200150 65480
rect 200350 65410 200360 65480
rect 200140 65360 200360 65410
rect 200640 65590 200860 65640
rect 200640 65520 200650 65590
rect 200850 65520 200860 65590
rect 200640 65480 200860 65520
rect 200640 65410 200650 65480
rect 200850 65410 200860 65480
rect 200640 65360 200860 65410
rect 201140 65590 201360 65640
rect 201140 65520 201150 65590
rect 201350 65520 201360 65590
rect 201140 65480 201360 65520
rect 201140 65410 201150 65480
rect 201350 65410 201360 65480
rect 201140 65360 201360 65410
rect 201640 65590 201860 65640
rect 201640 65520 201650 65590
rect 201850 65520 201860 65590
rect 201640 65480 201860 65520
rect 201640 65410 201650 65480
rect 201850 65410 201860 65480
rect 201640 65360 201860 65410
rect 202140 65590 202360 65640
rect 202140 65520 202150 65590
rect 202350 65520 202360 65590
rect 202140 65480 202360 65520
rect 202140 65410 202150 65480
rect 202350 65410 202360 65480
rect 202140 65360 202360 65410
rect 202640 65590 202860 65640
rect 202640 65520 202650 65590
rect 202850 65520 202860 65590
rect 202640 65480 202860 65520
rect 202640 65410 202650 65480
rect 202850 65410 202860 65480
rect 202640 65360 202860 65410
rect 203140 65590 203360 65640
rect 203140 65520 203150 65590
rect 203350 65520 203360 65590
rect 203140 65480 203360 65520
rect 203140 65410 203150 65480
rect 203350 65410 203360 65480
rect 203140 65360 203360 65410
rect 203640 65590 203860 65640
rect 203640 65520 203650 65590
rect 203850 65520 203860 65590
rect 203640 65480 203860 65520
rect 203640 65410 203650 65480
rect 203850 65410 203860 65480
rect 203640 65360 203860 65410
rect 204140 65590 204360 65640
rect 204140 65520 204150 65590
rect 204350 65520 204360 65590
rect 204140 65480 204360 65520
rect 204140 65410 204150 65480
rect 204350 65410 204360 65480
rect 204140 65360 204360 65410
rect 204640 65590 204860 65640
rect 204640 65520 204650 65590
rect 204850 65520 204860 65590
rect 204640 65480 204860 65520
rect 204640 65410 204650 65480
rect 204850 65410 204860 65480
rect 204640 65360 204860 65410
rect 205140 65590 205360 65640
rect 205140 65520 205150 65590
rect 205350 65520 205360 65590
rect 205140 65480 205360 65520
rect 205140 65410 205150 65480
rect 205350 65410 205360 65480
rect 205140 65360 205360 65410
rect 205640 65590 205860 65640
rect 205640 65520 205650 65590
rect 205850 65520 205860 65590
rect 205640 65480 205860 65520
rect 205640 65410 205650 65480
rect 205850 65410 205860 65480
rect 205640 65360 205860 65410
rect 206140 65590 206360 65640
rect 206140 65520 206150 65590
rect 206350 65520 206360 65590
rect 206140 65480 206360 65520
rect 206140 65410 206150 65480
rect 206350 65410 206360 65480
rect 206140 65360 206360 65410
rect 206640 65590 206860 65640
rect 206640 65520 206650 65590
rect 206850 65520 206860 65590
rect 206640 65480 206860 65520
rect 206640 65410 206650 65480
rect 206850 65410 206860 65480
rect 206640 65360 206860 65410
rect 207140 65590 207360 65640
rect 207140 65520 207150 65590
rect 207350 65520 207360 65590
rect 207140 65480 207360 65520
rect 207140 65410 207150 65480
rect 207350 65410 207360 65480
rect 207140 65360 207360 65410
rect 207640 65590 207860 65640
rect 207640 65520 207650 65590
rect 207850 65520 207860 65590
rect 207640 65480 207860 65520
rect 207640 65410 207650 65480
rect 207850 65410 207860 65480
rect 207640 65360 207860 65410
rect 190000 65350 208000 65360
rect 190000 65150 190020 65350
rect 190090 65150 190410 65350
rect 190480 65150 190520 65350
rect 190590 65150 190910 65350
rect 190980 65150 191020 65350
rect 191090 65150 191410 65350
rect 191480 65150 191520 65350
rect 191590 65150 191910 65350
rect 191980 65150 192020 65350
rect 192090 65150 192410 65350
rect 192480 65150 192520 65350
rect 192590 65150 192910 65350
rect 192980 65150 193020 65350
rect 193090 65150 193410 65350
rect 193480 65150 193520 65350
rect 193590 65150 193910 65350
rect 193980 65150 194020 65350
rect 194090 65150 194410 65350
rect 194480 65150 194520 65350
rect 194590 65150 194910 65350
rect 194980 65150 195020 65350
rect 195090 65150 195410 65350
rect 195480 65150 195520 65350
rect 195590 65150 195910 65350
rect 195980 65150 196020 65350
rect 196090 65150 196410 65350
rect 196480 65150 196520 65350
rect 196590 65150 196910 65350
rect 196980 65150 197020 65350
rect 197090 65150 197410 65350
rect 197480 65150 197520 65350
rect 197590 65150 197910 65350
rect 197980 65150 198020 65350
rect 198090 65150 198410 65350
rect 198480 65150 198520 65350
rect 198590 65150 198910 65350
rect 198980 65150 199020 65350
rect 199090 65150 199410 65350
rect 199480 65150 199520 65350
rect 199590 65150 199910 65350
rect 199980 65150 200020 65350
rect 200090 65150 200410 65350
rect 200480 65150 200520 65350
rect 200590 65150 200910 65350
rect 200980 65150 201020 65350
rect 201090 65150 201410 65350
rect 201480 65150 201520 65350
rect 201590 65150 201910 65350
rect 201980 65150 202020 65350
rect 202090 65150 202410 65350
rect 202480 65150 202520 65350
rect 202590 65150 202910 65350
rect 202980 65150 203020 65350
rect 203090 65150 203410 65350
rect 203480 65150 203520 65350
rect 203590 65150 203910 65350
rect 203980 65150 204020 65350
rect 204090 65150 204410 65350
rect 204480 65150 204520 65350
rect 204590 65150 204910 65350
rect 204980 65150 205020 65350
rect 205090 65150 205410 65350
rect 205480 65150 205520 65350
rect 205590 65150 205910 65350
rect 205980 65150 206020 65350
rect 206090 65150 206410 65350
rect 206480 65150 206520 65350
rect 206590 65150 206910 65350
rect 206980 65150 207020 65350
rect 207090 65150 207410 65350
rect 207480 65150 207520 65350
rect 207590 65150 207910 65350
rect 207980 65150 208000 65350
rect 190000 65140 208000 65150
rect 190140 65090 190360 65140
rect 190140 65020 190150 65090
rect 190350 65020 190360 65090
rect 190140 64980 190360 65020
rect 190140 64910 190150 64980
rect 190350 64910 190360 64980
rect 190140 64860 190360 64910
rect 190640 65090 190860 65140
rect 190640 65020 190650 65090
rect 190850 65020 190860 65090
rect 190640 64980 190860 65020
rect 190640 64910 190650 64980
rect 190850 64910 190860 64980
rect 190640 64860 190860 64910
rect 191140 65090 191360 65140
rect 191140 65020 191150 65090
rect 191350 65020 191360 65090
rect 191140 64980 191360 65020
rect 191140 64910 191150 64980
rect 191350 64910 191360 64980
rect 191140 64860 191360 64910
rect 191640 65090 191860 65140
rect 191640 65020 191650 65090
rect 191850 65020 191860 65090
rect 191640 64980 191860 65020
rect 191640 64910 191650 64980
rect 191850 64910 191860 64980
rect 191640 64860 191860 64910
rect 192140 65090 192360 65140
rect 192140 65020 192150 65090
rect 192350 65020 192360 65090
rect 192140 64980 192360 65020
rect 192140 64910 192150 64980
rect 192350 64910 192360 64980
rect 192140 64860 192360 64910
rect 192640 65090 192860 65140
rect 192640 65020 192650 65090
rect 192850 65020 192860 65090
rect 192640 64980 192860 65020
rect 192640 64910 192650 64980
rect 192850 64910 192860 64980
rect 192640 64860 192860 64910
rect 193140 65090 193360 65140
rect 193140 65020 193150 65090
rect 193350 65020 193360 65090
rect 193140 64980 193360 65020
rect 193140 64910 193150 64980
rect 193350 64910 193360 64980
rect 193140 64860 193360 64910
rect 193640 65090 193860 65140
rect 193640 65020 193650 65090
rect 193850 65020 193860 65090
rect 193640 64980 193860 65020
rect 193640 64910 193650 64980
rect 193850 64910 193860 64980
rect 193640 64860 193860 64910
rect 194140 65090 194360 65140
rect 194140 65020 194150 65090
rect 194350 65020 194360 65090
rect 194140 64980 194360 65020
rect 194140 64910 194150 64980
rect 194350 64910 194360 64980
rect 194140 64860 194360 64910
rect 194640 65090 194860 65140
rect 194640 65020 194650 65090
rect 194850 65020 194860 65090
rect 194640 64980 194860 65020
rect 194640 64910 194650 64980
rect 194850 64910 194860 64980
rect 194640 64860 194860 64910
rect 195140 65090 195360 65140
rect 195140 65020 195150 65090
rect 195350 65020 195360 65090
rect 195140 64980 195360 65020
rect 195140 64910 195150 64980
rect 195350 64910 195360 64980
rect 195140 64860 195360 64910
rect 195640 65090 195860 65140
rect 195640 65020 195650 65090
rect 195850 65020 195860 65090
rect 195640 64980 195860 65020
rect 195640 64910 195650 64980
rect 195850 64910 195860 64980
rect 195640 64860 195860 64910
rect 196140 65090 196360 65140
rect 196140 65020 196150 65090
rect 196350 65020 196360 65090
rect 196140 64980 196360 65020
rect 196140 64910 196150 64980
rect 196350 64910 196360 64980
rect 196140 64860 196360 64910
rect 196640 65090 196860 65140
rect 196640 65020 196650 65090
rect 196850 65020 196860 65090
rect 196640 64980 196860 65020
rect 196640 64910 196650 64980
rect 196850 64910 196860 64980
rect 196640 64860 196860 64910
rect 197140 65090 197360 65140
rect 197140 65020 197150 65090
rect 197350 65020 197360 65090
rect 197140 64980 197360 65020
rect 197140 64910 197150 64980
rect 197350 64910 197360 64980
rect 197140 64860 197360 64910
rect 197640 65090 197860 65140
rect 197640 65020 197650 65090
rect 197850 65020 197860 65090
rect 197640 64980 197860 65020
rect 197640 64910 197650 64980
rect 197850 64910 197860 64980
rect 197640 64860 197860 64910
rect 198140 65090 198360 65140
rect 198140 65020 198150 65090
rect 198350 65020 198360 65090
rect 198140 64980 198360 65020
rect 198140 64910 198150 64980
rect 198350 64910 198360 64980
rect 198140 64860 198360 64910
rect 198640 65090 198860 65140
rect 198640 65020 198650 65090
rect 198850 65020 198860 65090
rect 198640 64980 198860 65020
rect 198640 64910 198650 64980
rect 198850 64910 198860 64980
rect 198640 64860 198860 64910
rect 199140 65090 199360 65140
rect 199140 65020 199150 65090
rect 199350 65020 199360 65090
rect 199140 64980 199360 65020
rect 199140 64910 199150 64980
rect 199350 64910 199360 64980
rect 199140 64860 199360 64910
rect 199640 65090 199860 65140
rect 199640 65020 199650 65090
rect 199850 65020 199860 65090
rect 199640 64980 199860 65020
rect 199640 64910 199650 64980
rect 199850 64910 199860 64980
rect 199640 64860 199860 64910
rect 200140 65090 200360 65140
rect 200140 65020 200150 65090
rect 200350 65020 200360 65090
rect 200140 64980 200360 65020
rect 200140 64910 200150 64980
rect 200350 64910 200360 64980
rect 200140 64860 200360 64910
rect 200640 65090 200860 65140
rect 200640 65020 200650 65090
rect 200850 65020 200860 65090
rect 200640 64980 200860 65020
rect 200640 64910 200650 64980
rect 200850 64910 200860 64980
rect 200640 64860 200860 64910
rect 201140 65090 201360 65140
rect 201140 65020 201150 65090
rect 201350 65020 201360 65090
rect 201140 64980 201360 65020
rect 201140 64910 201150 64980
rect 201350 64910 201360 64980
rect 201140 64860 201360 64910
rect 201640 65090 201860 65140
rect 201640 65020 201650 65090
rect 201850 65020 201860 65090
rect 201640 64980 201860 65020
rect 201640 64910 201650 64980
rect 201850 64910 201860 64980
rect 201640 64860 201860 64910
rect 202140 65090 202360 65140
rect 202140 65020 202150 65090
rect 202350 65020 202360 65090
rect 202140 64980 202360 65020
rect 202140 64910 202150 64980
rect 202350 64910 202360 64980
rect 202140 64860 202360 64910
rect 202640 65090 202860 65140
rect 202640 65020 202650 65090
rect 202850 65020 202860 65090
rect 202640 64980 202860 65020
rect 202640 64910 202650 64980
rect 202850 64910 202860 64980
rect 202640 64860 202860 64910
rect 203140 65090 203360 65140
rect 203140 65020 203150 65090
rect 203350 65020 203360 65090
rect 203140 64980 203360 65020
rect 203140 64910 203150 64980
rect 203350 64910 203360 64980
rect 203140 64860 203360 64910
rect 203640 65090 203860 65140
rect 203640 65020 203650 65090
rect 203850 65020 203860 65090
rect 203640 64980 203860 65020
rect 203640 64910 203650 64980
rect 203850 64910 203860 64980
rect 203640 64860 203860 64910
rect 204140 65090 204360 65140
rect 204140 65020 204150 65090
rect 204350 65020 204360 65090
rect 204140 64980 204360 65020
rect 204140 64910 204150 64980
rect 204350 64910 204360 64980
rect 204140 64860 204360 64910
rect 204640 65090 204860 65140
rect 204640 65020 204650 65090
rect 204850 65020 204860 65090
rect 204640 64980 204860 65020
rect 204640 64910 204650 64980
rect 204850 64910 204860 64980
rect 204640 64860 204860 64910
rect 205140 65090 205360 65140
rect 205140 65020 205150 65090
rect 205350 65020 205360 65090
rect 205140 64980 205360 65020
rect 205140 64910 205150 64980
rect 205350 64910 205360 64980
rect 205140 64860 205360 64910
rect 205640 65090 205860 65140
rect 205640 65020 205650 65090
rect 205850 65020 205860 65090
rect 205640 64980 205860 65020
rect 205640 64910 205650 64980
rect 205850 64910 205860 64980
rect 205640 64860 205860 64910
rect 206140 65090 206360 65140
rect 206140 65020 206150 65090
rect 206350 65020 206360 65090
rect 206140 64980 206360 65020
rect 206140 64910 206150 64980
rect 206350 64910 206360 64980
rect 206140 64860 206360 64910
rect 206640 65090 206860 65140
rect 206640 65020 206650 65090
rect 206850 65020 206860 65090
rect 206640 64980 206860 65020
rect 206640 64910 206650 64980
rect 206850 64910 206860 64980
rect 206640 64860 206860 64910
rect 207140 65090 207360 65140
rect 207140 65020 207150 65090
rect 207350 65020 207360 65090
rect 207140 64980 207360 65020
rect 207140 64910 207150 64980
rect 207350 64910 207360 64980
rect 207140 64860 207360 64910
rect 207640 65090 207860 65140
rect 207640 65020 207650 65090
rect 207850 65020 207860 65090
rect 207640 64980 207860 65020
rect 207640 64910 207650 64980
rect 207850 64910 207860 64980
rect 207640 64860 207860 64910
rect 190000 64850 208000 64860
rect 190000 64650 190020 64850
rect 190090 64650 190410 64850
rect 190480 64650 190520 64850
rect 190590 64650 190910 64850
rect 190980 64650 191020 64850
rect 191090 64650 191410 64850
rect 191480 64650 191520 64850
rect 191590 64650 191910 64850
rect 191980 64650 192020 64850
rect 192090 64650 192410 64850
rect 192480 64650 192520 64850
rect 192590 64650 192910 64850
rect 192980 64650 193020 64850
rect 193090 64650 193410 64850
rect 193480 64650 193520 64850
rect 193590 64650 193910 64850
rect 193980 64650 194020 64850
rect 194090 64650 194410 64850
rect 194480 64650 194520 64850
rect 194590 64650 194910 64850
rect 194980 64650 195020 64850
rect 195090 64650 195410 64850
rect 195480 64650 195520 64850
rect 195590 64650 195910 64850
rect 195980 64650 196020 64850
rect 196090 64650 196410 64850
rect 196480 64650 196520 64850
rect 196590 64650 196910 64850
rect 196980 64650 197020 64850
rect 197090 64650 197410 64850
rect 197480 64650 197520 64850
rect 197590 64650 197910 64850
rect 197980 64650 198020 64850
rect 198090 64650 198410 64850
rect 198480 64650 198520 64850
rect 198590 64650 198910 64850
rect 198980 64650 199020 64850
rect 199090 64650 199410 64850
rect 199480 64650 199520 64850
rect 199590 64650 199910 64850
rect 199980 64650 200020 64850
rect 200090 64650 200410 64850
rect 200480 64650 200520 64850
rect 200590 64650 200910 64850
rect 200980 64650 201020 64850
rect 201090 64650 201410 64850
rect 201480 64650 201520 64850
rect 201590 64650 201910 64850
rect 201980 64650 202020 64850
rect 202090 64650 202410 64850
rect 202480 64650 202520 64850
rect 202590 64650 202910 64850
rect 202980 64650 203020 64850
rect 203090 64650 203410 64850
rect 203480 64650 203520 64850
rect 203590 64650 203910 64850
rect 203980 64650 204020 64850
rect 204090 64650 204410 64850
rect 204480 64650 204520 64850
rect 204590 64650 204910 64850
rect 204980 64650 205020 64850
rect 205090 64650 205410 64850
rect 205480 64650 205520 64850
rect 205590 64650 205910 64850
rect 205980 64650 206020 64850
rect 206090 64650 206410 64850
rect 206480 64650 206520 64850
rect 206590 64650 206910 64850
rect 206980 64650 207020 64850
rect 207090 64650 207410 64850
rect 207480 64650 207520 64850
rect 207590 64650 207910 64850
rect 207980 64650 208000 64850
rect 190000 64640 208000 64650
rect 190140 64590 190360 64640
rect 190140 64520 190150 64590
rect 190350 64520 190360 64590
rect 190140 64480 190360 64520
rect 190140 64410 190150 64480
rect 190350 64410 190360 64480
rect 190140 64360 190360 64410
rect 190640 64590 190860 64640
rect 190640 64520 190650 64590
rect 190850 64520 190860 64590
rect 190640 64480 190860 64520
rect 190640 64410 190650 64480
rect 190850 64410 190860 64480
rect 190640 64360 190860 64410
rect 191140 64590 191360 64640
rect 191140 64520 191150 64590
rect 191350 64520 191360 64590
rect 191140 64480 191360 64520
rect 191140 64410 191150 64480
rect 191350 64410 191360 64480
rect 191140 64360 191360 64410
rect 191640 64590 191860 64640
rect 191640 64520 191650 64590
rect 191850 64520 191860 64590
rect 191640 64480 191860 64520
rect 191640 64410 191650 64480
rect 191850 64410 191860 64480
rect 191640 64360 191860 64410
rect 192140 64590 192360 64640
rect 192140 64520 192150 64590
rect 192350 64520 192360 64590
rect 192140 64480 192360 64520
rect 192140 64410 192150 64480
rect 192350 64410 192360 64480
rect 192140 64360 192360 64410
rect 192640 64590 192860 64640
rect 192640 64520 192650 64590
rect 192850 64520 192860 64590
rect 192640 64480 192860 64520
rect 192640 64410 192650 64480
rect 192850 64410 192860 64480
rect 192640 64360 192860 64410
rect 193140 64590 193360 64640
rect 193140 64520 193150 64590
rect 193350 64520 193360 64590
rect 193140 64480 193360 64520
rect 193140 64410 193150 64480
rect 193350 64410 193360 64480
rect 193140 64360 193360 64410
rect 193640 64590 193860 64640
rect 193640 64520 193650 64590
rect 193850 64520 193860 64590
rect 193640 64480 193860 64520
rect 193640 64410 193650 64480
rect 193850 64410 193860 64480
rect 193640 64360 193860 64410
rect 194140 64590 194360 64640
rect 194140 64520 194150 64590
rect 194350 64520 194360 64590
rect 194140 64480 194360 64520
rect 194140 64410 194150 64480
rect 194350 64410 194360 64480
rect 194140 64360 194360 64410
rect 194640 64590 194860 64640
rect 194640 64520 194650 64590
rect 194850 64520 194860 64590
rect 194640 64480 194860 64520
rect 194640 64410 194650 64480
rect 194850 64410 194860 64480
rect 194640 64360 194860 64410
rect 195140 64590 195360 64640
rect 195140 64520 195150 64590
rect 195350 64520 195360 64590
rect 195140 64480 195360 64520
rect 195140 64410 195150 64480
rect 195350 64410 195360 64480
rect 195140 64360 195360 64410
rect 195640 64590 195860 64640
rect 195640 64520 195650 64590
rect 195850 64520 195860 64590
rect 195640 64480 195860 64520
rect 195640 64410 195650 64480
rect 195850 64410 195860 64480
rect 195640 64360 195860 64410
rect 196140 64590 196360 64640
rect 196140 64520 196150 64590
rect 196350 64520 196360 64590
rect 196140 64480 196360 64520
rect 196140 64410 196150 64480
rect 196350 64410 196360 64480
rect 196140 64360 196360 64410
rect 196640 64590 196860 64640
rect 196640 64520 196650 64590
rect 196850 64520 196860 64590
rect 196640 64480 196860 64520
rect 196640 64410 196650 64480
rect 196850 64410 196860 64480
rect 196640 64360 196860 64410
rect 197140 64590 197360 64640
rect 197140 64520 197150 64590
rect 197350 64520 197360 64590
rect 197140 64480 197360 64520
rect 197140 64410 197150 64480
rect 197350 64410 197360 64480
rect 197140 64360 197360 64410
rect 197640 64590 197860 64640
rect 197640 64520 197650 64590
rect 197850 64520 197860 64590
rect 197640 64480 197860 64520
rect 197640 64410 197650 64480
rect 197850 64410 197860 64480
rect 197640 64360 197860 64410
rect 198140 64590 198360 64640
rect 198140 64520 198150 64590
rect 198350 64520 198360 64590
rect 198140 64480 198360 64520
rect 198140 64410 198150 64480
rect 198350 64410 198360 64480
rect 198140 64360 198360 64410
rect 198640 64590 198860 64640
rect 198640 64520 198650 64590
rect 198850 64520 198860 64590
rect 198640 64480 198860 64520
rect 198640 64410 198650 64480
rect 198850 64410 198860 64480
rect 198640 64360 198860 64410
rect 199140 64590 199360 64640
rect 199140 64520 199150 64590
rect 199350 64520 199360 64590
rect 199140 64480 199360 64520
rect 199140 64410 199150 64480
rect 199350 64410 199360 64480
rect 199140 64360 199360 64410
rect 199640 64590 199860 64640
rect 199640 64520 199650 64590
rect 199850 64520 199860 64590
rect 199640 64480 199860 64520
rect 199640 64410 199650 64480
rect 199850 64410 199860 64480
rect 199640 64360 199860 64410
rect 200140 64590 200360 64640
rect 200140 64520 200150 64590
rect 200350 64520 200360 64590
rect 200140 64480 200360 64520
rect 200140 64410 200150 64480
rect 200350 64410 200360 64480
rect 200140 64360 200360 64410
rect 200640 64590 200860 64640
rect 200640 64520 200650 64590
rect 200850 64520 200860 64590
rect 200640 64480 200860 64520
rect 200640 64410 200650 64480
rect 200850 64410 200860 64480
rect 200640 64360 200860 64410
rect 201140 64590 201360 64640
rect 201140 64520 201150 64590
rect 201350 64520 201360 64590
rect 201140 64480 201360 64520
rect 201140 64410 201150 64480
rect 201350 64410 201360 64480
rect 201140 64360 201360 64410
rect 201640 64590 201860 64640
rect 201640 64520 201650 64590
rect 201850 64520 201860 64590
rect 201640 64480 201860 64520
rect 201640 64410 201650 64480
rect 201850 64410 201860 64480
rect 201640 64360 201860 64410
rect 202140 64590 202360 64640
rect 202140 64520 202150 64590
rect 202350 64520 202360 64590
rect 202140 64480 202360 64520
rect 202140 64410 202150 64480
rect 202350 64410 202360 64480
rect 202140 64360 202360 64410
rect 202640 64590 202860 64640
rect 202640 64520 202650 64590
rect 202850 64520 202860 64590
rect 202640 64480 202860 64520
rect 202640 64410 202650 64480
rect 202850 64410 202860 64480
rect 202640 64360 202860 64410
rect 203140 64590 203360 64640
rect 203140 64520 203150 64590
rect 203350 64520 203360 64590
rect 203140 64480 203360 64520
rect 203140 64410 203150 64480
rect 203350 64410 203360 64480
rect 203140 64360 203360 64410
rect 203640 64590 203860 64640
rect 203640 64520 203650 64590
rect 203850 64520 203860 64590
rect 203640 64480 203860 64520
rect 203640 64410 203650 64480
rect 203850 64410 203860 64480
rect 203640 64360 203860 64410
rect 204140 64590 204360 64640
rect 204140 64520 204150 64590
rect 204350 64520 204360 64590
rect 204140 64480 204360 64520
rect 204140 64410 204150 64480
rect 204350 64410 204360 64480
rect 204140 64360 204360 64410
rect 204640 64590 204860 64640
rect 204640 64520 204650 64590
rect 204850 64520 204860 64590
rect 204640 64480 204860 64520
rect 204640 64410 204650 64480
rect 204850 64410 204860 64480
rect 204640 64360 204860 64410
rect 205140 64590 205360 64640
rect 205140 64520 205150 64590
rect 205350 64520 205360 64590
rect 205140 64480 205360 64520
rect 205140 64410 205150 64480
rect 205350 64410 205360 64480
rect 205140 64360 205360 64410
rect 205640 64590 205860 64640
rect 205640 64520 205650 64590
rect 205850 64520 205860 64590
rect 205640 64480 205860 64520
rect 205640 64410 205650 64480
rect 205850 64410 205860 64480
rect 205640 64360 205860 64410
rect 206140 64590 206360 64640
rect 206140 64520 206150 64590
rect 206350 64520 206360 64590
rect 206140 64480 206360 64520
rect 206140 64410 206150 64480
rect 206350 64410 206360 64480
rect 206140 64360 206360 64410
rect 206640 64590 206860 64640
rect 206640 64520 206650 64590
rect 206850 64520 206860 64590
rect 206640 64480 206860 64520
rect 206640 64410 206650 64480
rect 206850 64410 206860 64480
rect 206640 64360 206860 64410
rect 207140 64590 207360 64640
rect 207140 64520 207150 64590
rect 207350 64520 207360 64590
rect 207140 64480 207360 64520
rect 207140 64410 207150 64480
rect 207350 64410 207360 64480
rect 207140 64360 207360 64410
rect 207640 64590 207860 64640
rect 207640 64520 207650 64590
rect 207850 64520 207860 64590
rect 207640 64480 207860 64520
rect 207640 64410 207650 64480
rect 207850 64410 207860 64480
rect 207640 64360 207860 64410
rect 190000 64350 208000 64360
rect 190000 64150 190020 64350
rect 190090 64150 190410 64350
rect 190480 64150 190520 64350
rect 190590 64150 190910 64350
rect 190980 64150 191020 64350
rect 191090 64150 191410 64350
rect 191480 64150 191520 64350
rect 191590 64150 191910 64350
rect 191980 64150 192020 64350
rect 192090 64150 192410 64350
rect 192480 64150 192520 64350
rect 192590 64150 192910 64350
rect 192980 64150 193020 64350
rect 193090 64150 193410 64350
rect 193480 64150 193520 64350
rect 193590 64150 193910 64350
rect 193980 64150 194020 64350
rect 194090 64150 194410 64350
rect 194480 64150 194520 64350
rect 194590 64150 194910 64350
rect 194980 64150 195020 64350
rect 195090 64150 195410 64350
rect 195480 64150 195520 64350
rect 195590 64150 195910 64350
rect 195980 64150 196020 64350
rect 196090 64150 196410 64350
rect 196480 64150 196520 64350
rect 196590 64150 196910 64350
rect 196980 64150 197020 64350
rect 197090 64150 197410 64350
rect 197480 64150 197520 64350
rect 197590 64150 197910 64350
rect 197980 64150 198020 64350
rect 198090 64150 198410 64350
rect 198480 64150 198520 64350
rect 198590 64150 198910 64350
rect 198980 64150 199020 64350
rect 199090 64150 199410 64350
rect 199480 64150 199520 64350
rect 199590 64150 199910 64350
rect 199980 64150 200020 64350
rect 200090 64150 200410 64350
rect 200480 64150 200520 64350
rect 200590 64150 200910 64350
rect 200980 64150 201020 64350
rect 201090 64150 201410 64350
rect 201480 64150 201520 64350
rect 201590 64150 201910 64350
rect 201980 64150 202020 64350
rect 202090 64150 202410 64350
rect 202480 64150 202520 64350
rect 202590 64150 202910 64350
rect 202980 64150 203020 64350
rect 203090 64150 203410 64350
rect 203480 64150 203520 64350
rect 203590 64150 203910 64350
rect 203980 64150 204020 64350
rect 204090 64150 204410 64350
rect 204480 64150 204520 64350
rect 204590 64150 204910 64350
rect 204980 64150 205020 64350
rect 205090 64150 205410 64350
rect 205480 64150 205520 64350
rect 205590 64150 205910 64350
rect 205980 64150 206020 64350
rect 206090 64150 206410 64350
rect 206480 64150 206520 64350
rect 206590 64150 206910 64350
rect 206980 64150 207020 64350
rect 207090 64150 207410 64350
rect 207480 64150 207520 64350
rect 207590 64150 207910 64350
rect 207980 64150 208000 64350
rect 190000 64140 208000 64150
rect 190140 64090 190360 64140
rect 190140 64020 190150 64090
rect 190350 64020 190360 64090
rect 190140 64000 190360 64020
rect 190640 64090 190860 64140
rect 190640 64020 190650 64090
rect 190850 64020 190860 64090
rect 190640 64000 190860 64020
rect 191140 64090 191360 64140
rect 191140 64020 191150 64090
rect 191350 64020 191360 64090
rect 191140 64000 191360 64020
rect 191640 64090 191860 64140
rect 191640 64020 191650 64090
rect 191850 64020 191860 64090
rect 191640 64000 191860 64020
rect 192140 64090 192360 64140
rect 192140 64020 192150 64090
rect 192350 64020 192360 64090
rect 192140 64000 192360 64020
rect 192640 64090 192860 64140
rect 192640 64020 192650 64090
rect 192850 64020 192860 64090
rect 192640 64000 192860 64020
rect 193140 64090 193360 64140
rect 193140 64020 193150 64090
rect 193350 64020 193360 64090
rect 193140 64000 193360 64020
rect 193640 64090 193860 64140
rect 193640 64020 193650 64090
rect 193850 64020 193860 64090
rect 193640 64000 193860 64020
rect 194140 64090 194360 64140
rect 194140 64020 194150 64090
rect 194350 64020 194360 64090
rect 194140 64000 194360 64020
rect 194640 64090 194860 64140
rect 194640 64020 194650 64090
rect 194850 64020 194860 64090
rect 194640 64000 194860 64020
rect 195140 64090 195360 64140
rect 195140 64020 195150 64090
rect 195350 64020 195360 64090
rect 195140 64000 195360 64020
rect 195640 64090 195860 64140
rect 195640 64020 195650 64090
rect 195850 64020 195860 64090
rect 195640 64000 195860 64020
rect 196140 64090 196360 64140
rect 196140 64020 196150 64090
rect 196350 64020 196360 64090
rect 196140 64000 196360 64020
rect 196640 64090 196860 64140
rect 196640 64020 196650 64090
rect 196850 64020 196860 64090
rect 196640 64000 196860 64020
rect 197140 64090 197360 64140
rect 197140 64020 197150 64090
rect 197350 64020 197360 64090
rect 197140 64000 197360 64020
rect 197640 64090 197860 64140
rect 197640 64020 197650 64090
rect 197850 64020 197860 64090
rect 197640 64000 197860 64020
rect 198140 64090 198360 64140
rect 198140 64020 198150 64090
rect 198350 64020 198360 64090
rect 198140 64000 198360 64020
rect 198640 64090 198860 64140
rect 198640 64020 198650 64090
rect 198850 64020 198860 64090
rect 198640 64000 198860 64020
rect 199140 64090 199360 64140
rect 199140 64020 199150 64090
rect 199350 64020 199360 64090
rect 199140 64000 199360 64020
rect 199640 64090 199860 64140
rect 199640 64020 199650 64090
rect 199850 64020 199860 64090
rect 199640 64000 199860 64020
rect 200140 64090 200360 64140
rect 200140 64020 200150 64090
rect 200350 64020 200360 64090
rect 200140 64000 200360 64020
rect 200640 64090 200860 64140
rect 200640 64020 200650 64090
rect 200850 64020 200860 64090
rect 200640 64000 200860 64020
rect 201140 64090 201360 64140
rect 201140 64020 201150 64090
rect 201350 64020 201360 64090
rect 201140 64000 201360 64020
rect 201640 64090 201860 64140
rect 201640 64020 201650 64090
rect 201850 64020 201860 64090
rect 201640 64000 201860 64020
rect 202140 64090 202360 64140
rect 202140 64020 202150 64090
rect 202350 64020 202360 64090
rect 202140 64000 202360 64020
rect 202640 64090 202860 64140
rect 202640 64020 202650 64090
rect 202850 64020 202860 64090
rect 202640 64000 202860 64020
rect 203140 64090 203360 64140
rect 203140 64020 203150 64090
rect 203350 64020 203360 64090
rect 203140 64000 203360 64020
rect 203640 64090 203860 64140
rect 203640 64020 203650 64090
rect 203850 64020 203860 64090
rect 203640 64000 203860 64020
rect 204140 64090 204360 64140
rect 204140 64020 204150 64090
rect 204350 64020 204360 64090
rect 204140 63980 204360 64020
rect 204140 63910 204150 63980
rect 204350 63910 204360 63980
rect 204140 63860 204360 63910
rect 204640 64090 204860 64140
rect 204640 64020 204650 64090
rect 204850 64020 204860 64090
rect 204640 63980 204860 64020
rect 204640 63910 204650 63980
rect 204850 63910 204860 63980
rect 204640 63860 204860 63910
rect 205140 64090 205360 64140
rect 205140 64020 205150 64090
rect 205350 64020 205360 64090
rect 205140 63980 205360 64020
rect 205140 63910 205150 63980
rect 205350 63910 205360 63980
rect 205140 63860 205360 63910
rect 205640 64090 205860 64140
rect 205640 64020 205650 64090
rect 205850 64020 205860 64090
rect 205640 63980 205860 64020
rect 205640 63910 205650 63980
rect 205850 63910 205860 63980
rect 205640 63860 205860 63910
rect 206140 64090 206360 64140
rect 206140 64020 206150 64090
rect 206350 64020 206360 64090
rect 206140 63980 206360 64020
rect 206140 63910 206150 63980
rect 206350 63910 206360 63980
rect 206140 63860 206360 63910
rect 206640 64090 206860 64140
rect 206640 64020 206650 64090
rect 206850 64020 206860 64090
rect 206640 63980 206860 64020
rect 206640 63910 206650 63980
rect 206850 63910 206860 63980
rect 206640 63860 206860 63910
rect 207140 64090 207360 64140
rect 207140 64020 207150 64090
rect 207350 64020 207360 64090
rect 207140 63980 207360 64020
rect 207140 63910 207150 63980
rect 207350 63910 207360 63980
rect 207140 63860 207360 63910
rect 207640 64090 207860 64140
rect 207640 64020 207650 64090
rect 207850 64020 207860 64090
rect 207640 63980 207860 64020
rect 207640 63910 207650 63980
rect 207850 63910 207860 63980
rect 207640 63860 207860 63910
rect 204000 63850 208000 63860
rect 204000 63650 204020 63850
rect 204090 63650 204410 63850
rect 204480 63650 204520 63850
rect 204590 63650 204910 63850
rect 204980 63650 205020 63850
rect 205090 63650 205410 63850
rect 205480 63650 205520 63850
rect 205590 63650 205910 63850
rect 205980 63650 206020 63850
rect 206090 63650 206410 63850
rect 206480 63650 206520 63850
rect 206590 63650 206910 63850
rect 206980 63650 207020 63850
rect 207090 63650 207410 63850
rect 207480 63650 207520 63850
rect 207590 63650 207910 63850
rect 207980 63650 208000 63850
rect 204000 63640 208000 63650
rect 204140 63590 204360 63640
rect 204140 63520 204150 63590
rect 204350 63520 204360 63590
rect 204140 63480 204360 63520
rect 204140 63410 204150 63480
rect 204350 63410 204360 63480
rect 204140 63360 204360 63410
rect 204640 63590 204860 63640
rect 204640 63520 204650 63590
rect 204850 63520 204860 63590
rect 204640 63480 204860 63520
rect 204640 63410 204650 63480
rect 204850 63410 204860 63480
rect 204640 63360 204860 63410
rect 205140 63590 205360 63640
rect 205140 63520 205150 63590
rect 205350 63520 205360 63590
rect 205140 63480 205360 63520
rect 205140 63410 205150 63480
rect 205350 63410 205360 63480
rect 205140 63360 205360 63410
rect 205640 63590 205860 63640
rect 205640 63520 205650 63590
rect 205850 63520 205860 63590
rect 205640 63480 205860 63520
rect 205640 63410 205650 63480
rect 205850 63410 205860 63480
rect 205640 63360 205860 63410
rect 206140 63590 206360 63640
rect 206140 63520 206150 63590
rect 206350 63520 206360 63590
rect 206140 63480 206360 63520
rect 206140 63410 206150 63480
rect 206350 63410 206360 63480
rect 206140 63360 206360 63410
rect 206640 63590 206860 63640
rect 206640 63520 206650 63590
rect 206850 63520 206860 63590
rect 206640 63480 206860 63520
rect 206640 63410 206650 63480
rect 206850 63410 206860 63480
rect 206640 63360 206860 63410
rect 207140 63590 207360 63640
rect 207140 63520 207150 63590
rect 207350 63520 207360 63590
rect 207140 63480 207360 63520
rect 207140 63410 207150 63480
rect 207350 63410 207360 63480
rect 207140 63360 207360 63410
rect 207640 63590 207860 63640
rect 207640 63520 207650 63590
rect 207850 63520 207860 63590
rect 207640 63480 207860 63520
rect 207640 63410 207650 63480
rect 207850 63410 207860 63480
rect 207640 63360 207860 63410
rect 204000 63350 208000 63360
rect 204000 63150 204020 63350
rect 204090 63150 204410 63350
rect 204480 63150 204520 63350
rect 204590 63150 204910 63350
rect 204980 63150 205020 63350
rect 205090 63150 205410 63350
rect 205480 63150 205520 63350
rect 205590 63150 205910 63350
rect 205980 63150 206020 63350
rect 206090 63150 206410 63350
rect 206480 63150 206520 63350
rect 206590 63150 206910 63350
rect 206980 63150 207020 63350
rect 207090 63150 207410 63350
rect 207480 63150 207520 63350
rect 207590 63150 207910 63350
rect 207980 63150 208000 63350
rect 204000 63140 208000 63150
rect 204140 63090 204360 63140
rect 204140 63020 204150 63090
rect 204350 63020 204360 63090
rect 204140 62980 204360 63020
rect 204140 62910 204150 62980
rect 204350 62910 204360 62980
rect 204140 62860 204360 62910
rect 204640 63090 204860 63140
rect 204640 63020 204650 63090
rect 204850 63020 204860 63090
rect 204640 62980 204860 63020
rect 204640 62910 204650 62980
rect 204850 62910 204860 62980
rect 204640 62860 204860 62910
rect 205140 63090 205360 63140
rect 205140 63020 205150 63090
rect 205350 63020 205360 63090
rect 205140 62980 205360 63020
rect 205140 62910 205150 62980
rect 205350 62910 205360 62980
rect 205140 62860 205360 62910
rect 205640 63090 205860 63140
rect 205640 63020 205650 63090
rect 205850 63020 205860 63090
rect 205640 62980 205860 63020
rect 205640 62910 205650 62980
rect 205850 62910 205860 62980
rect 205640 62860 205860 62910
rect 206140 63090 206360 63140
rect 206140 63020 206150 63090
rect 206350 63020 206360 63090
rect 206140 62980 206360 63020
rect 206140 62910 206150 62980
rect 206350 62910 206360 62980
rect 206140 62860 206360 62910
rect 206640 63090 206860 63140
rect 206640 63020 206650 63090
rect 206850 63020 206860 63090
rect 206640 62980 206860 63020
rect 206640 62910 206650 62980
rect 206850 62910 206860 62980
rect 206640 62860 206860 62910
rect 207140 63090 207360 63140
rect 207140 63020 207150 63090
rect 207350 63020 207360 63090
rect 207140 62980 207360 63020
rect 207140 62910 207150 62980
rect 207350 62910 207360 62980
rect 207140 62860 207360 62910
rect 207640 63090 207860 63140
rect 207640 63020 207650 63090
rect 207850 63020 207860 63090
rect 207640 62980 207860 63020
rect 207640 62910 207650 62980
rect 207850 62910 207860 62980
rect 207640 62860 207860 62910
rect 204000 62850 208000 62860
rect 204000 62650 204020 62850
rect 204090 62650 204410 62850
rect 204480 62650 204520 62850
rect 204590 62650 204910 62850
rect 204980 62650 205020 62850
rect 205090 62650 205410 62850
rect 205480 62650 205520 62850
rect 205590 62650 205910 62850
rect 205980 62650 206020 62850
rect 206090 62650 206410 62850
rect 206480 62650 206520 62850
rect 206590 62650 206910 62850
rect 206980 62650 207020 62850
rect 207090 62650 207410 62850
rect 207480 62650 207520 62850
rect 207590 62650 207910 62850
rect 207980 62650 208000 62850
rect 204000 62640 208000 62650
rect 204140 62590 204360 62640
rect 204140 62520 204150 62590
rect 204350 62520 204360 62590
rect 204140 62480 204360 62520
rect 204140 62410 204150 62480
rect 204350 62410 204360 62480
rect 204140 62360 204360 62410
rect 204640 62590 204860 62640
rect 204640 62520 204650 62590
rect 204850 62520 204860 62590
rect 204640 62480 204860 62520
rect 204640 62410 204650 62480
rect 204850 62410 204860 62480
rect 204640 62360 204860 62410
rect 205140 62590 205360 62640
rect 205140 62520 205150 62590
rect 205350 62520 205360 62590
rect 205140 62480 205360 62520
rect 205140 62410 205150 62480
rect 205350 62410 205360 62480
rect 205140 62360 205360 62410
rect 205640 62590 205860 62640
rect 205640 62520 205650 62590
rect 205850 62520 205860 62590
rect 205640 62480 205860 62520
rect 205640 62410 205650 62480
rect 205850 62410 205860 62480
rect 205640 62360 205860 62410
rect 206140 62590 206360 62640
rect 206140 62520 206150 62590
rect 206350 62520 206360 62590
rect 206140 62480 206360 62520
rect 206140 62410 206150 62480
rect 206350 62410 206360 62480
rect 206140 62360 206360 62410
rect 206640 62590 206860 62640
rect 206640 62520 206650 62590
rect 206850 62520 206860 62590
rect 206640 62480 206860 62520
rect 206640 62410 206650 62480
rect 206850 62410 206860 62480
rect 206640 62360 206860 62410
rect 207140 62590 207360 62640
rect 207140 62520 207150 62590
rect 207350 62520 207360 62590
rect 207140 62480 207360 62520
rect 207140 62410 207150 62480
rect 207350 62410 207360 62480
rect 207140 62360 207360 62410
rect 207640 62590 207860 62640
rect 207640 62520 207650 62590
rect 207850 62520 207860 62590
rect 207640 62480 207860 62520
rect 207640 62410 207650 62480
rect 207850 62410 207860 62480
rect 207640 62360 207860 62410
rect 204000 62350 208000 62360
rect 204000 62150 204020 62350
rect 204090 62150 204410 62350
rect 204480 62150 204520 62350
rect 204590 62150 204910 62350
rect 204980 62150 205020 62350
rect 205090 62150 205410 62350
rect 205480 62150 205520 62350
rect 205590 62150 205910 62350
rect 205980 62150 206020 62350
rect 206090 62150 206410 62350
rect 206480 62150 206520 62350
rect 206590 62150 206910 62350
rect 206980 62150 207020 62350
rect 207090 62150 207410 62350
rect 207480 62150 207520 62350
rect 207590 62150 207910 62350
rect 207980 62150 208000 62350
rect 204000 62140 208000 62150
rect 204140 62090 204360 62140
rect 204140 62020 204150 62090
rect 204350 62020 204360 62090
rect 204140 61980 204360 62020
rect 204140 61910 204150 61980
rect 204350 61910 204360 61980
rect 204140 61860 204360 61910
rect 204640 62090 204860 62140
rect 204640 62020 204650 62090
rect 204850 62020 204860 62090
rect 204640 61980 204860 62020
rect 204640 61910 204650 61980
rect 204850 61910 204860 61980
rect 204640 61860 204860 61910
rect 205140 62090 205360 62140
rect 205140 62020 205150 62090
rect 205350 62020 205360 62090
rect 205140 61980 205360 62020
rect 205140 61910 205150 61980
rect 205350 61910 205360 61980
rect 205140 61860 205360 61910
rect 205640 62090 205860 62140
rect 205640 62020 205650 62090
rect 205850 62020 205860 62090
rect 205640 61980 205860 62020
rect 205640 61910 205650 61980
rect 205850 61910 205860 61980
rect 205640 61860 205860 61910
rect 206140 62090 206360 62140
rect 206140 62020 206150 62090
rect 206350 62020 206360 62090
rect 206140 61980 206360 62020
rect 206140 61910 206150 61980
rect 206350 61910 206360 61980
rect 206140 61860 206360 61910
rect 206640 62090 206860 62140
rect 206640 62020 206650 62090
rect 206850 62020 206860 62090
rect 206640 61980 206860 62020
rect 206640 61910 206650 61980
rect 206850 61910 206860 61980
rect 206640 61860 206860 61910
rect 207140 62090 207360 62140
rect 207140 62020 207150 62090
rect 207350 62020 207360 62090
rect 207140 61980 207360 62020
rect 207140 61910 207150 61980
rect 207350 61910 207360 61980
rect 207140 61860 207360 61910
rect 207640 62090 207860 62140
rect 207640 62020 207650 62090
rect 207850 62020 207860 62090
rect 207640 61980 207860 62020
rect 207640 61910 207650 61980
rect 207850 61910 207860 61980
rect 207640 61860 207860 61910
rect 204000 61850 208000 61860
rect 204000 61650 204020 61850
rect 204090 61650 204410 61850
rect 204480 61650 204520 61850
rect 204590 61650 204910 61850
rect 204980 61650 205020 61850
rect 205090 61650 205410 61850
rect 205480 61650 205520 61850
rect 205590 61650 205910 61850
rect 205980 61650 206020 61850
rect 206090 61650 206410 61850
rect 206480 61650 206520 61850
rect 206590 61650 206910 61850
rect 206980 61650 207020 61850
rect 207090 61650 207410 61850
rect 207480 61650 207520 61850
rect 207590 61650 207910 61850
rect 207980 61650 208000 61850
rect 204000 61640 208000 61650
rect 204140 61590 204360 61640
rect 204140 61520 204150 61590
rect 204350 61520 204360 61590
rect 204140 61480 204360 61520
rect 204140 61410 204150 61480
rect 204350 61410 204360 61480
rect 204140 61360 204360 61410
rect 204640 61590 204860 61640
rect 204640 61520 204650 61590
rect 204850 61520 204860 61590
rect 204640 61480 204860 61520
rect 204640 61410 204650 61480
rect 204850 61410 204860 61480
rect 204640 61360 204860 61410
rect 205140 61590 205360 61640
rect 205140 61520 205150 61590
rect 205350 61520 205360 61590
rect 205140 61480 205360 61520
rect 205140 61410 205150 61480
rect 205350 61410 205360 61480
rect 205140 61360 205360 61410
rect 205640 61590 205860 61640
rect 205640 61520 205650 61590
rect 205850 61520 205860 61590
rect 205640 61480 205860 61520
rect 205640 61410 205650 61480
rect 205850 61410 205860 61480
rect 205640 61360 205860 61410
rect 206140 61590 206360 61640
rect 206140 61520 206150 61590
rect 206350 61520 206360 61590
rect 206140 61480 206360 61520
rect 206140 61410 206150 61480
rect 206350 61410 206360 61480
rect 206140 61360 206360 61410
rect 206640 61590 206860 61640
rect 206640 61520 206650 61590
rect 206850 61520 206860 61590
rect 206640 61480 206860 61520
rect 206640 61410 206650 61480
rect 206850 61410 206860 61480
rect 206640 61360 206860 61410
rect 207140 61590 207360 61640
rect 207140 61520 207150 61590
rect 207350 61520 207360 61590
rect 207140 61480 207360 61520
rect 207140 61410 207150 61480
rect 207350 61410 207360 61480
rect 207140 61360 207360 61410
rect 207640 61590 207860 61640
rect 207640 61520 207650 61590
rect 207850 61520 207860 61590
rect 207640 61480 207860 61520
rect 207640 61410 207650 61480
rect 207850 61410 207860 61480
rect 207640 61360 207860 61410
rect 204000 61350 208000 61360
rect 204000 61150 204020 61350
rect 204090 61150 204410 61350
rect 204480 61150 204520 61350
rect 204590 61150 204910 61350
rect 204980 61150 205020 61350
rect 205090 61150 205410 61350
rect 205480 61150 205520 61350
rect 205590 61150 205910 61350
rect 205980 61150 206020 61350
rect 206090 61150 206410 61350
rect 206480 61150 206520 61350
rect 206590 61150 206910 61350
rect 206980 61150 207020 61350
rect 207090 61150 207410 61350
rect 207480 61150 207520 61350
rect 207590 61150 207910 61350
rect 207980 61150 208000 61350
rect 204000 61140 208000 61150
rect 204140 61090 204360 61140
rect 204140 61020 204150 61090
rect 204350 61020 204360 61090
rect 204140 60980 204360 61020
rect 204140 60910 204150 60980
rect 204350 60910 204360 60980
rect 204140 60860 204360 60910
rect 204640 61090 204860 61140
rect 204640 61020 204650 61090
rect 204850 61020 204860 61090
rect 204640 60980 204860 61020
rect 204640 60910 204650 60980
rect 204850 60910 204860 60980
rect 204640 60860 204860 60910
rect 205140 61090 205360 61140
rect 205140 61020 205150 61090
rect 205350 61020 205360 61090
rect 205140 60980 205360 61020
rect 205140 60910 205150 60980
rect 205350 60910 205360 60980
rect 205140 60860 205360 60910
rect 205640 61090 205860 61140
rect 205640 61020 205650 61090
rect 205850 61020 205860 61090
rect 205640 60980 205860 61020
rect 205640 60910 205650 60980
rect 205850 60910 205860 60980
rect 205640 60860 205860 60910
rect 206140 61090 206360 61140
rect 206140 61020 206150 61090
rect 206350 61020 206360 61090
rect 206140 60980 206360 61020
rect 206140 60910 206150 60980
rect 206350 60910 206360 60980
rect 206140 60860 206360 60910
rect 206640 61090 206860 61140
rect 206640 61020 206650 61090
rect 206850 61020 206860 61090
rect 206640 60980 206860 61020
rect 206640 60910 206650 60980
rect 206850 60910 206860 60980
rect 206640 60860 206860 60910
rect 207140 61090 207360 61140
rect 207140 61020 207150 61090
rect 207350 61020 207360 61090
rect 207140 60980 207360 61020
rect 207140 60910 207150 60980
rect 207350 60910 207360 60980
rect 207140 60860 207360 60910
rect 207640 61090 207860 61140
rect 207640 61020 207650 61090
rect 207850 61020 207860 61090
rect 207640 60980 207860 61020
rect 207640 60910 207650 60980
rect 207850 60910 207860 60980
rect 207640 60860 207860 60910
rect 204000 60850 208000 60860
rect 204000 60650 204020 60850
rect 204090 60650 204410 60850
rect 204480 60650 204520 60850
rect 204590 60650 204910 60850
rect 204980 60650 205020 60850
rect 205090 60650 205410 60850
rect 205480 60650 205520 60850
rect 205590 60650 205910 60850
rect 205980 60650 206020 60850
rect 206090 60650 206410 60850
rect 206480 60650 206520 60850
rect 206590 60650 206910 60850
rect 206980 60650 207020 60850
rect 207090 60650 207410 60850
rect 207480 60650 207520 60850
rect 207590 60650 207910 60850
rect 207980 60650 208000 60850
rect 204000 60640 208000 60650
rect 204140 60590 204360 60640
rect 204140 60520 204150 60590
rect 204350 60520 204360 60590
rect 204140 60480 204360 60520
rect 204140 60410 204150 60480
rect 204350 60410 204360 60480
rect 204140 60360 204360 60410
rect 204640 60590 204860 60640
rect 204640 60520 204650 60590
rect 204850 60520 204860 60590
rect 204640 60480 204860 60520
rect 204640 60410 204650 60480
rect 204850 60410 204860 60480
rect 204640 60360 204860 60410
rect 205140 60590 205360 60640
rect 205140 60520 205150 60590
rect 205350 60520 205360 60590
rect 205140 60480 205360 60520
rect 205140 60410 205150 60480
rect 205350 60410 205360 60480
rect 205140 60360 205360 60410
rect 205640 60590 205860 60640
rect 205640 60520 205650 60590
rect 205850 60520 205860 60590
rect 205640 60480 205860 60520
rect 205640 60410 205650 60480
rect 205850 60410 205860 60480
rect 205640 60360 205860 60410
rect 206140 60590 206360 60640
rect 206140 60520 206150 60590
rect 206350 60520 206360 60590
rect 206140 60480 206360 60520
rect 206140 60410 206150 60480
rect 206350 60410 206360 60480
rect 206140 60360 206360 60410
rect 206640 60590 206860 60640
rect 206640 60520 206650 60590
rect 206850 60520 206860 60590
rect 206640 60480 206860 60520
rect 206640 60410 206650 60480
rect 206850 60410 206860 60480
rect 206640 60360 206860 60410
rect 207140 60590 207360 60640
rect 207140 60520 207150 60590
rect 207350 60520 207360 60590
rect 207140 60480 207360 60520
rect 207140 60410 207150 60480
rect 207350 60410 207360 60480
rect 207140 60360 207360 60410
rect 207640 60590 207860 60640
rect 207640 60520 207650 60590
rect 207850 60520 207860 60590
rect 207640 60480 207860 60520
rect 207640 60410 207650 60480
rect 207850 60410 207860 60480
rect 207640 60360 207860 60410
rect 204000 60350 208000 60360
rect 204000 60150 204020 60350
rect 204090 60150 204410 60350
rect 204480 60150 204520 60350
rect 204590 60150 204910 60350
rect 204980 60150 205020 60350
rect 205090 60150 205410 60350
rect 205480 60150 205520 60350
rect 205590 60150 205910 60350
rect 205980 60150 206020 60350
rect 206090 60150 206410 60350
rect 206480 60150 206520 60350
rect 206590 60150 206910 60350
rect 206980 60150 207020 60350
rect 207090 60150 207410 60350
rect 207480 60150 207520 60350
rect 207590 60150 207910 60350
rect 207980 60150 208000 60350
rect 204000 60140 208000 60150
rect 204140 60090 204360 60140
rect 204140 60020 204150 60090
rect 204350 60020 204360 60090
rect 204140 59980 204360 60020
rect 204140 59910 204150 59980
rect 204350 59910 204360 59980
rect 204140 59860 204360 59910
rect 204640 60090 204860 60140
rect 204640 60020 204650 60090
rect 204850 60020 204860 60090
rect 204640 59980 204860 60020
rect 204640 59910 204650 59980
rect 204850 59910 204860 59980
rect 204640 59860 204860 59910
rect 205140 60090 205360 60140
rect 205140 60020 205150 60090
rect 205350 60020 205360 60090
rect 205140 59980 205360 60020
rect 205140 59910 205150 59980
rect 205350 59910 205360 59980
rect 205140 59860 205360 59910
rect 205640 60090 205860 60140
rect 205640 60020 205650 60090
rect 205850 60020 205860 60090
rect 205640 59980 205860 60020
rect 205640 59910 205650 59980
rect 205850 59910 205860 59980
rect 205640 59860 205860 59910
rect 206140 60090 206360 60140
rect 206140 60020 206150 60090
rect 206350 60020 206360 60090
rect 206140 59980 206360 60020
rect 206140 59910 206150 59980
rect 206350 59910 206360 59980
rect 206140 59860 206360 59910
rect 206640 60090 206860 60140
rect 206640 60020 206650 60090
rect 206850 60020 206860 60090
rect 206640 59980 206860 60020
rect 206640 59910 206650 59980
rect 206850 59910 206860 59980
rect 206640 59860 206860 59910
rect 207140 60090 207360 60140
rect 207140 60020 207150 60090
rect 207350 60020 207360 60090
rect 207140 59980 207360 60020
rect 207140 59910 207150 59980
rect 207350 59910 207360 59980
rect 207140 59860 207360 59910
rect 207640 60090 207860 60140
rect 207640 60020 207650 60090
rect 207850 60020 207860 60090
rect 207640 59980 207860 60020
rect 207640 59910 207650 59980
rect 207850 59910 207860 59980
rect 207640 59860 207860 59910
rect 204000 59850 208000 59860
rect 204000 59650 204020 59850
rect 204090 59650 204410 59850
rect 204480 59650 204520 59850
rect 204590 59650 204910 59850
rect 204980 59650 205020 59850
rect 205090 59650 205410 59850
rect 205480 59650 205520 59850
rect 205590 59650 205910 59850
rect 205980 59650 206020 59850
rect 206090 59650 206410 59850
rect 206480 59650 206520 59850
rect 206590 59650 206910 59850
rect 206980 59650 207020 59850
rect 207090 59650 207410 59850
rect 207480 59650 207520 59850
rect 207590 59650 207910 59850
rect 207980 59650 208000 59850
rect 204000 59640 208000 59650
rect 204140 59590 204360 59640
rect 204140 59520 204150 59590
rect 204350 59520 204360 59590
rect 204140 59480 204360 59520
rect 204140 59410 204150 59480
rect 204350 59410 204360 59480
rect 204140 59360 204360 59410
rect 204640 59590 204860 59640
rect 204640 59520 204650 59590
rect 204850 59520 204860 59590
rect 204640 59480 204860 59520
rect 204640 59410 204650 59480
rect 204850 59410 204860 59480
rect 204640 59360 204860 59410
rect 205140 59590 205360 59640
rect 205140 59520 205150 59590
rect 205350 59520 205360 59590
rect 205140 59480 205360 59520
rect 205140 59410 205150 59480
rect 205350 59410 205360 59480
rect 205140 59360 205360 59410
rect 205640 59590 205860 59640
rect 205640 59520 205650 59590
rect 205850 59520 205860 59590
rect 205640 59480 205860 59520
rect 205640 59410 205650 59480
rect 205850 59410 205860 59480
rect 205640 59360 205860 59410
rect 206140 59590 206360 59640
rect 206140 59520 206150 59590
rect 206350 59520 206360 59590
rect 206140 59480 206360 59520
rect 206140 59410 206150 59480
rect 206350 59410 206360 59480
rect 206140 59360 206360 59410
rect 206640 59590 206860 59640
rect 206640 59520 206650 59590
rect 206850 59520 206860 59590
rect 206640 59480 206860 59520
rect 206640 59410 206650 59480
rect 206850 59410 206860 59480
rect 206640 59360 206860 59410
rect 207140 59590 207360 59640
rect 207140 59520 207150 59590
rect 207350 59520 207360 59590
rect 207140 59480 207360 59520
rect 207140 59410 207150 59480
rect 207350 59410 207360 59480
rect 207140 59360 207360 59410
rect 207640 59590 207860 59640
rect 207640 59520 207650 59590
rect 207850 59520 207860 59590
rect 207640 59480 207860 59520
rect 207640 59410 207650 59480
rect 207850 59410 207860 59480
rect 207640 59360 207860 59410
rect 204000 59350 208000 59360
rect 204000 59150 204020 59350
rect 204090 59150 204410 59350
rect 204480 59150 204520 59350
rect 204590 59150 204910 59350
rect 204980 59150 205020 59350
rect 205090 59150 205410 59350
rect 205480 59150 205520 59350
rect 205590 59150 205910 59350
rect 205980 59150 206020 59350
rect 206090 59150 206410 59350
rect 206480 59150 206520 59350
rect 206590 59150 206910 59350
rect 206980 59150 207020 59350
rect 207090 59150 207410 59350
rect 207480 59150 207520 59350
rect 207590 59150 207910 59350
rect 207980 59150 208000 59350
rect 204000 59140 208000 59150
rect 204140 59090 204360 59140
rect 204140 59020 204150 59090
rect 204350 59020 204360 59090
rect 204140 58980 204360 59020
rect 204140 58910 204150 58980
rect 204350 58910 204360 58980
rect 204140 58860 204360 58910
rect 204640 59090 204860 59140
rect 204640 59020 204650 59090
rect 204850 59020 204860 59090
rect 204640 58980 204860 59020
rect 204640 58910 204650 58980
rect 204850 58910 204860 58980
rect 204640 58860 204860 58910
rect 205140 59090 205360 59140
rect 205140 59020 205150 59090
rect 205350 59020 205360 59090
rect 205140 58980 205360 59020
rect 205140 58910 205150 58980
rect 205350 58910 205360 58980
rect 205140 58860 205360 58910
rect 205640 59090 205860 59140
rect 205640 59020 205650 59090
rect 205850 59020 205860 59090
rect 205640 58980 205860 59020
rect 205640 58910 205650 58980
rect 205850 58910 205860 58980
rect 205640 58860 205860 58910
rect 206140 59090 206360 59140
rect 206140 59020 206150 59090
rect 206350 59020 206360 59090
rect 206140 58980 206360 59020
rect 206140 58910 206150 58980
rect 206350 58910 206360 58980
rect 206140 58860 206360 58910
rect 206640 59090 206860 59140
rect 206640 59020 206650 59090
rect 206850 59020 206860 59090
rect 206640 58980 206860 59020
rect 206640 58910 206650 58980
rect 206850 58910 206860 58980
rect 206640 58860 206860 58910
rect 207140 59090 207360 59140
rect 207140 59020 207150 59090
rect 207350 59020 207360 59090
rect 207140 58980 207360 59020
rect 207140 58910 207150 58980
rect 207350 58910 207360 58980
rect 207140 58860 207360 58910
rect 207640 59090 207860 59140
rect 207640 59020 207650 59090
rect 207850 59020 207860 59090
rect 207640 58980 207860 59020
rect 207640 58910 207650 58980
rect 207850 58910 207860 58980
rect 207640 58860 207860 58910
rect 204000 58850 208000 58860
rect 204000 58650 204020 58850
rect 204090 58650 204410 58850
rect 204480 58650 204520 58850
rect 204590 58650 204910 58850
rect 204980 58650 205020 58850
rect 205090 58650 205410 58850
rect 205480 58650 205520 58850
rect 205590 58650 205910 58850
rect 205980 58650 206020 58850
rect 206090 58650 206410 58850
rect 206480 58650 206520 58850
rect 206590 58650 206910 58850
rect 206980 58650 207020 58850
rect 207090 58650 207410 58850
rect 207480 58650 207520 58850
rect 207590 58650 207910 58850
rect 207980 58650 208000 58850
rect 204000 58640 208000 58650
rect 204140 58590 204360 58640
rect 204140 58520 204150 58590
rect 204350 58520 204360 58590
rect 204140 58480 204360 58520
rect 204140 58410 204150 58480
rect 204350 58410 204360 58480
rect 204140 58360 204360 58410
rect 204640 58590 204860 58640
rect 204640 58520 204650 58590
rect 204850 58520 204860 58590
rect 204640 58480 204860 58520
rect 204640 58410 204650 58480
rect 204850 58410 204860 58480
rect 204640 58360 204860 58410
rect 205140 58590 205360 58640
rect 205140 58520 205150 58590
rect 205350 58520 205360 58590
rect 205140 58480 205360 58520
rect 205140 58410 205150 58480
rect 205350 58410 205360 58480
rect 205140 58360 205360 58410
rect 205640 58590 205860 58640
rect 205640 58520 205650 58590
rect 205850 58520 205860 58590
rect 205640 58480 205860 58520
rect 205640 58410 205650 58480
rect 205850 58410 205860 58480
rect 205640 58360 205860 58410
rect 206140 58590 206360 58640
rect 206140 58520 206150 58590
rect 206350 58520 206360 58590
rect 206140 58480 206360 58520
rect 206140 58410 206150 58480
rect 206350 58410 206360 58480
rect 206140 58360 206360 58410
rect 206640 58590 206860 58640
rect 206640 58520 206650 58590
rect 206850 58520 206860 58590
rect 206640 58480 206860 58520
rect 206640 58410 206650 58480
rect 206850 58410 206860 58480
rect 206640 58360 206860 58410
rect 207140 58590 207360 58640
rect 207140 58520 207150 58590
rect 207350 58520 207360 58590
rect 207140 58480 207360 58520
rect 207140 58410 207150 58480
rect 207350 58410 207360 58480
rect 207140 58360 207360 58410
rect 207640 58590 207860 58640
rect 207640 58520 207650 58590
rect 207850 58520 207860 58590
rect 207640 58480 207860 58520
rect 207640 58410 207650 58480
rect 207850 58410 207860 58480
rect 207640 58360 207860 58410
rect 204000 58350 208000 58360
rect 204000 58150 204020 58350
rect 204090 58150 204410 58350
rect 204480 58150 204520 58350
rect 204590 58150 204910 58350
rect 204980 58150 205020 58350
rect 205090 58150 205410 58350
rect 205480 58150 205520 58350
rect 205590 58150 205910 58350
rect 205980 58150 206020 58350
rect 206090 58150 206410 58350
rect 206480 58150 206520 58350
rect 206590 58150 206910 58350
rect 206980 58150 207020 58350
rect 207090 58150 207410 58350
rect 207480 58150 207520 58350
rect 207590 58150 207910 58350
rect 207980 58150 208000 58350
rect 204000 58140 208000 58150
rect 204140 58090 204360 58140
rect 204140 58020 204150 58090
rect 204350 58020 204360 58090
rect 204140 57980 204360 58020
rect 204140 57910 204150 57980
rect 204350 57910 204360 57980
rect 204140 57860 204360 57910
rect 204640 58090 204860 58140
rect 204640 58020 204650 58090
rect 204850 58020 204860 58090
rect 204640 57980 204860 58020
rect 204640 57910 204650 57980
rect 204850 57910 204860 57980
rect 204640 57860 204860 57910
rect 205140 58090 205360 58140
rect 205140 58020 205150 58090
rect 205350 58020 205360 58090
rect 205140 57980 205360 58020
rect 205140 57910 205150 57980
rect 205350 57910 205360 57980
rect 205140 57860 205360 57910
rect 205640 58090 205860 58140
rect 205640 58020 205650 58090
rect 205850 58020 205860 58090
rect 205640 57980 205860 58020
rect 205640 57910 205650 57980
rect 205850 57910 205860 57980
rect 205640 57860 205860 57910
rect 206140 58090 206360 58140
rect 206140 58020 206150 58090
rect 206350 58020 206360 58090
rect 206140 57980 206360 58020
rect 206140 57910 206150 57980
rect 206350 57910 206360 57980
rect 206140 57860 206360 57910
rect 206640 58090 206860 58140
rect 206640 58020 206650 58090
rect 206850 58020 206860 58090
rect 206640 57980 206860 58020
rect 206640 57910 206650 57980
rect 206850 57910 206860 57980
rect 206640 57860 206860 57910
rect 207140 58090 207360 58140
rect 207140 58020 207150 58090
rect 207350 58020 207360 58090
rect 207140 57980 207360 58020
rect 207140 57910 207150 57980
rect 207350 57910 207360 57980
rect 207140 57860 207360 57910
rect 207640 58090 207860 58140
rect 207640 58020 207650 58090
rect 207850 58020 207860 58090
rect 207640 57980 207860 58020
rect 207640 57910 207650 57980
rect 207850 57910 207860 57980
rect 207640 57860 207860 57910
rect 204000 57850 208000 57860
rect 204000 57650 204020 57850
rect 204090 57650 204410 57850
rect 204480 57650 204520 57850
rect 204590 57650 204910 57850
rect 204980 57650 205020 57850
rect 205090 57650 205410 57850
rect 205480 57650 205520 57850
rect 205590 57650 205910 57850
rect 205980 57650 206020 57850
rect 206090 57650 206410 57850
rect 206480 57650 206520 57850
rect 206590 57650 206910 57850
rect 206980 57650 207020 57850
rect 207090 57650 207410 57850
rect 207480 57650 207520 57850
rect 207590 57650 207910 57850
rect 207980 57650 208000 57850
rect 204000 57640 208000 57650
rect 204140 57590 204360 57640
rect 204140 57520 204150 57590
rect 204350 57520 204360 57590
rect 204140 57480 204360 57520
rect 204140 57410 204150 57480
rect 204350 57410 204360 57480
rect 204140 57360 204360 57410
rect 204640 57590 204860 57640
rect 204640 57520 204650 57590
rect 204850 57520 204860 57590
rect 204640 57480 204860 57520
rect 204640 57410 204650 57480
rect 204850 57410 204860 57480
rect 204640 57360 204860 57410
rect 205140 57590 205360 57640
rect 205140 57520 205150 57590
rect 205350 57520 205360 57590
rect 205140 57480 205360 57520
rect 205140 57410 205150 57480
rect 205350 57410 205360 57480
rect 205140 57360 205360 57410
rect 205640 57590 205860 57640
rect 205640 57520 205650 57590
rect 205850 57520 205860 57590
rect 205640 57480 205860 57520
rect 205640 57410 205650 57480
rect 205850 57410 205860 57480
rect 205640 57360 205860 57410
rect 206140 57590 206360 57640
rect 206140 57520 206150 57590
rect 206350 57520 206360 57590
rect 206140 57480 206360 57520
rect 206140 57410 206150 57480
rect 206350 57410 206360 57480
rect 206140 57360 206360 57410
rect 206640 57590 206860 57640
rect 206640 57520 206650 57590
rect 206850 57520 206860 57590
rect 206640 57480 206860 57520
rect 206640 57410 206650 57480
rect 206850 57410 206860 57480
rect 206640 57360 206860 57410
rect 207140 57590 207360 57640
rect 207140 57520 207150 57590
rect 207350 57520 207360 57590
rect 207140 57480 207360 57520
rect 207140 57410 207150 57480
rect 207350 57410 207360 57480
rect 207140 57360 207360 57410
rect 207640 57590 207860 57640
rect 207640 57520 207650 57590
rect 207850 57520 207860 57590
rect 207640 57480 207860 57520
rect 207640 57410 207650 57480
rect 207850 57410 207860 57480
rect 207640 57360 207860 57410
rect 204000 57350 208000 57360
rect 204000 57150 204020 57350
rect 204090 57150 204410 57350
rect 204480 57150 204520 57350
rect 204590 57150 204910 57350
rect 204980 57150 205020 57350
rect 205090 57150 205410 57350
rect 205480 57150 205520 57350
rect 205590 57150 205910 57350
rect 205980 57150 206020 57350
rect 206090 57150 206410 57350
rect 206480 57150 206520 57350
rect 206590 57150 206910 57350
rect 206980 57150 207020 57350
rect 207090 57150 207410 57350
rect 207480 57150 207520 57350
rect 207590 57150 207910 57350
rect 207980 57150 208000 57350
rect 204000 57140 208000 57150
rect 204140 57090 204360 57140
rect 204140 57020 204150 57090
rect 204350 57020 204360 57090
rect 204140 56980 204360 57020
rect 204140 56910 204150 56980
rect 204350 56910 204360 56980
rect 204140 56860 204360 56910
rect 204640 57090 204860 57140
rect 204640 57020 204650 57090
rect 204850 57020 204860 57090
rect 204640 56980 204860 57020
rect 204640 56910 204650 56980
rect 204850 56910 204860 56980
rect 204640 56860 204860 56910
rect 205140 57090 205360 57140
rect 205140 57020 205150 57090
rect 205350 57020 205360 57090
rect 205140 56980 205360 57020
rect 205140 56910 205150 56980
rect 205350 56910 205360 56980
rect 205140 56860 205360 56910
rect 205640 57090 205860 57140
rect 205640 57020 205650 57090
rect 205850 57020 205860 57090
rect 205640 56980 205860 57020
rect 205640 56910 205650 56980
rect 205850 56910 205860 56980
rect 205640 56860 205860 56910
rect 206140 57090 206360 57140
rect 206140 57020 206150 57090
rect 206350 57020 206360 57090
rect 206140 56980 206360 57020
rect 206140 56910 206150 56980
rect 206350 56910 206360 56980
rect 206140 56860 206360 56910
rect 206640 57090 206860 57140
rect 206640 57020 206650 57090
rect 206850 57020 206860 57090
rect 206640 56980 206860 57020
rect 206640 56910 206650 56980
rect 206850 56910 206860 56980
rect 206640 56860 206860 56910
rect 207140 57090 207360 57140
rect 207140 57020 207150 57090
rect 207350 57020 207360 57090
rect 207140 56980 207360 57020
rect 207140 56910 207150 56980
rect 207350 56910 207360 56980
rect 207140 56860 207360 56910
rect 207640 57090 207860 57140
rect 207640 57020 207650 57090
rect 207850 57020 207860 57090
rect 207640 56980 207860 57020
rect 207640 56910 207650 56980
rect 207850 56910 207860 56980
rect 207640 56860 207860 56910
rect 204000 56850 208000 56860
rect 204000 56650 204020 56850
rect 204090 56650 204410 56850
rect 204480 56650 204520 56850
rect 204590 56650 204910 56850
rect 204980 56650 205020 56850
rect 205090 56650 205410 56850
rect 205480 56650 205520 56850
rect 205590 56650 205910 56850
rect 205980 56650 206020 56850
rect 206090 56650 206410 56850
rect 206480 56650 206520 56850
rect 206590 56650 206910 56850
rect 206980 56650 207020 56850
rect 207090 56650 207410 56850
rect 207480 56650 207520 56850
rect 207590 56650 207910 56850
rect 207980 56650 208000 56850
rect 204000 56640 208000 56650
rect 204140 56590 204360 56640
rect 204140 56520 204150 56590
rect 204350 56520 204360 56590
rect 204140 56480 204360 56520
rect 204140 56410 204150 56480
rect 204350 56410 204360 56480
rect 204140 56360 204360 56410
rect 204640 56590 204860 56640
rect 204640 56520 204650 56590
rect 204850 56520 204860 56590
rect 204640 56480 204860 56520
rect 204640 56410 204650 56480
rect 204850 56410 204860 56480
rect 204640 56360 204860 56410
rect 205140 56590 205360 56640
rect 205140 56520 205150 56590
rect 205350 56520 205360 56590
rect 205140 56480 205360 56520
rect 205140 56410 205150 56480
rect 205350 56410 205360 56480
rect 205140 56360 205360 56410
rect 205640 56590 205860 56640
rect 205640 56520 205650 56590
rect 205850 56520 205860 56590
rect 205640 56480 205860 56520
rect 205640 56410 205650 56480
rect 205850 56410 205860 56480
rect 205640 56360 205860 56410
rect 206140 56590 206360 56640
rect 206140 56520 206150 56590
rect 206350 56520 206360 56590
rect 206140 56480 206360 56520
rect 206140 56410 206150 56480
rect 206350 56410 206360 56480
rect 206140 56360 206360 56410
rect 206640 56590 206860 56640
rect 206640 56520 206650 56590
rect 206850 56520 206860 56590
rect 206640 56480 206860 56520
rect 206640 56410 206650 56480
rect 206850 56410 206860 56480
rect 206640 56360 206860 56410
rect 207140 56590 207360 56640
rect 207140 56520 207150 56590
rect 207350 56520 207360 56590
rect 207140 56480 207360 56520
rect 207140 56410 207150 56480
rect 207350 56410 207360 56480
rect 207140 56360 207360 56410
rect 207640 56590 207860 56640
rect 207640 56520 207650 56590
rect 207850 56520 207860 56590
rect 207640 56480 207860 56520
rect 207640 56410 207650 56480
rect 207850 56410 207860 56480
rect 207640 56360 207860 56410
rect 204000 56350 208000 56360
rect 204000 56150 204020 56350
rect 204090 56150 204410 56350
rect 204480 56150 204520 56350
rect 204590 56150 204910 56350
rect 204980 56150 205020 56350
rect 205090 56150 205410 56350
rect 205480 56150 205520 56350
rect 205590 56150 205910 56350
rect 205980 56150 206020 56350
rect 206090 56150 206410 56350
rect 206480 56150 206520 56350
rect 206590 56150 206910 56350
rect 206980 56150 207020 56350
rect 207090 56150 207410 56350
rect 207480 56150 207520 56350
rect 207590 56150 207910 56350
rect 207980 56150 208000 56350
rect 204000 56140 208000 56150
rect 204140 56090 204360 56140
rect 204140 56020 204150 56090
rect 204350 56020 204360 56090
rect 204140 55980 204360 56020
rect 204140 55910 204150 55980
rect 204350 55910 204360 55980
rect 204140 55860 204360 55910
rect 204640 56090 204860 56140
rect 204640 56020 204650 56090
rect 204850 56020 204860 56090
rect 204640 55980 204860 56020
rect 204640 55910 204650 55980
rect 204850 55910 204860 55980
rect 204640 55860 204860 55910
rect 205140 56090 205360 56140
rect 205140 56020 205150 56090
rect 205350 56020 205360 56090
rect 205140 55980 205360 56020
rect 205140 55910 205150 55980
rect 205350 55910 205360 55980
rect 205140 55860 205360 55910
rect 205640 56090 205860 56140
rect 205640 56020 205650 56090
rect 205850 56020 205860 56090
rect 205640 55980 205860 56020
rect 205640 55910 205650 55980
rect 205850 55910 205860 55980
rect 205640 55860 205860 55910
rect 206140 56090 206360 56140
rect 206140 56020 206150 56090
rect 206350 56020 206360 56090
rect 206140 55980 206360 56020
rect 206140 55910 206150 55980
rect 206350 55910 206360 55980
rect 206140 55860 206360 55910
rect 206640 56090 206860 56140
rect 206640 56020 206650 56090
rect 206850 56020 206860 56090
rect 206640 55980 206860 56020
rect 206640 55910 206650 55980
rect 206850 55910 206860 55980
rect 206640 55860 206860 55910
rect 207140 56090 207360 56140
rect 207140 56020 207150 56090
rect 207350 56020 207360 56090
rect 207140 55980 207360 56020
rect 207140 55910 207150 55980
rect 207350 55910 207360 55980
rect 207140 55860 207360 55910
rect 207640 56090 207860 56140
rect 207640 56020 207650 56090
rect 207850 56020 207860 56090
rect 207640 55980 207860 56020
rect 207640 55910 207650 55980
rect 207850 55910 207860 55980
rect 207640 55860 207860 55910
rect 204000 55850 208000 55860
rect 204000 55650 204020 55850
rect 204090 55650 204410 55850
rect 204480 55650 204520 55850
rect 204590 55650 204910 55850
rect 204980 55650 205020 55850
rect 205090 55650 205410 55850
rect 205480 55650 205520 55850
rect 205590 55650 205910 55850
rect 205980 55650 206020 55850
rect 206090 55650 206410 55850
rect 206480 55650 206520 55850
rect 206590 55650 206910 55850
rect 206980 55650 207020 55850
rect 207090 55650 207410 55850
rect 207480 55650 207520 55850
rect 207590 55650 207910 55850
rect 207980 55650 208000 55850
rect 204000 55640 208000 55650
rect 204140 55590 204360 55640
rect 204140 55520 204150 55590
rect 204350 55520 204360 55590
rect 204140 55480 204360 55520
rect 204140 55410 204150 55480
rect 204350 55410 204360 55480
rect 204140 55360 204360 55410
rect 204640 55590 204860 55640
rect 204640 55520 204650 55590
rect 204850 55520 204860 55590
rect 204640 55480 204860 55520
rect 204640 55410 204650 55480
rect 204850 55410 204860 55480
rect 204640 55360 204860 55410
rect 205140 55590 205360 55640
rect 205140 55520 205150 55590
rect 205350 55520 205360 55590
rect 205140 55480 205360 55520
rect 205140 55410 205150 55480
rect 205350 55410 205360 55480
rect 205140 55360 205360 55410
rect 205640 55590 205860 55640
rect 205640 55520 205650 55590
rect 205850 55520 205860 55590
rect 205640 55480 205860 55520
rect 205640 55410 205650 55480
rect 205850 55410 205860 55480
rect 205640 55360 205860 55410
rect 206140 55590 206360 55640
rect 206140 55520 206150 55590
rect 206350 55520 206360 55590
rect 206140 55480 206360 55520
rect 206140 55410 206150 55480
rect 206350 55410 206360 55480
rect 206140 55360 206360 55410
rect 206640 55590 206860 55640
rect 206640 55520 206650 55590
rect 206850 55520 206860 55590
rect 206640 55480 206860 55520
rect 206640 55410 206650 55480
rect 206850 55410 206860 55480
rect 206640 55360 206860 55410
rect 207140 55590 207360 55640
rect 207140 55520 207150 55590
rect 207350 55520 207360 55590
rect 207140 55480 207360 55520
rect 207140 55410 207150 55480
rect 207350 55410 207360 55480
rect 207140 55360 207360 55410
rect 207640 55590 207860 55640
rect 207640 55520 207650 55590
rect 207850 55520 207860 55590
rect 207640 55480 207860 55520
rect 207640 55410 207650 55480
rect 207850 55410 207860 55480
rect 207640 55360 207860 55410
rect 204000 55350 208000 55360
rect 204000 55150 204020 55350
rect 204090 55150 204410 55350
rect 204480 55150 204520 55350
rect 204590 55150 204910 55350
rect 204980 55150 205020 55350
rect 205090 55150 205410 55350
rect 205480 55150 205520 55350
rect 205590 55150 205910 55350
rect 205980 55150 206020 55350
rect 206090 55150 206410 55350
rect 206480 55150 206520 55350
rect 206590 55150 206910 55350
rect 206980 55150 207020 55350
rect 207090 55150 207410 55350
rect 207480 55150 207520 55350
rect 207590 55150 207910 55350
rect 207980 55150 208000 55350
rect 204000 55140 208000 55150
rect 204140 55090 204360 55140
rect 204140 55020 204150 55090
rect 204350 55020 204360 55090
rect 204140 54980 204360 55020
rect 204140 54910 204150 54980
rect 204350 54910 204360 54980
rect 204140 54860 204360 54910
rect 204640 55090 204860 55140
rect 204640 55020 204650 55090
rect 204850 55020 204860 55090
rect 204640 54980 204860 55020
rect 204640 54910 204650 54980
rect 204850 54910 204860 54980
rect 204640 54860 204860 54910
rect 205140 55090 205360 55140
rect 205140 55020 205150 55090
rect 205350 55020 205360 55090
rect 205140 54980 205360 55020
rect 205140 54910 205150 54980
rect 205350 54910 205360 54980
rect 205140 54860 205360 54910
rect 205640 55090 205860 55140
rect 205640 55020 205650 55090
rect 205850 55020 205860 55090
rect 205640 54980 205860 55020
rect 205640 54910 205650 54980
rect 205850 54910 205860 54980
rect 205640 54860 205860 54910
rect 206140 55090 206360 55140
rect 206140 55020 206150 55090
rect 206350 55020 206360 55090
rect 206140 54980 206360 55020
rect 206140 54910 206150 54980
rect 206350 54910 206360 54980
rect 206140 54860 206360 54910
rect 206640 55090 206860 55140
rect 206640 55020 206650 55090
rect 206850 55020 206860 55090
rect 206640 54980 206860 55020
rect 206640 54910 206650 54980
rect 206850 54910 206860 54980
rect 206640 54860 206860 54910
rect 207140 55090 207360 55140
rect 207140 55020 207150 55090
rect 207350 55020 207360 55090
rect 207140 54980 207360 55020
rect 207140 54910 207150 54980
rect 207350 54910 207360 54980
rect 207140 54860 207360 54910
rect 207640 55090 207860 55140
rect 207640 55020 207650 55090
rect 207850 55020 207860 55090
rect 207640 54980 207860 55020
rect 207640 54910 207650 54980
rect 207850 54910 207860 54980
rect 207640 54860 207860 54910
rect 204000 54850 208000 54860
rect 204000 54650 204020 54850
rect 204090 54650 204410 54850
rect 204480 54650 204520 54850
rect 204590 54650 204910 54850
rect 204980 54650 205020 54850
rect 205090 54650 205410 54850
rect 205480 54650 205520 54850
rect 205590 54650 205910 54850
rect 205980 54650 206020 54850
rect 206090 54650 206410 54850
rect 206480 54650 206520 54850
rect 206590 54650 206910 54850
rect 206980 54650 207020 54850
rect 207090 54650 207410 54850
rect 207480 54650 207520 54850
rect 207590 54650 207910 54850
rect 207980 54650 208000 54850
rect 204000 54640 208000 54650
rect 204140 54590 204360 54640
rect 204140 54520 204150 54590
rect 204350 54520 204360 54590
rect 204140 54480 204360 54520
rect 204140 54410 204150 54480
rect 204350 54410 204360 54480
rect 204140 54360 204360 54410
rect 204640 54590 204860 54640
rect 204640 54520 204650 54590
rect 204850 54520 204860 54590
rect 204640 54480 204860 54520
rect 204640 54410 204650 54480
rect 204850 54410 204860 54480
rect 204640 54360 204860 54410
rect 205140 54590 205360 54640
rect 205140 54520 205150 54590
rect 205350 54520 205360 54590
rect 205140 54480 205360 54520
rect 205140 54410 205150 54480
rect 205350 54410 205360 54480
rect 205140 54360 205360 54410
rect 205640 54590 205860 54640
rect 205640 54520 205650 54590
rect 205850 54520 205860 54590
rect 205640 54480 205860 54520
rect 205640 54410 205650 54480
rect 205850 54410 205860 54480
rect 205640 54360 205860 54410
rect 206140 54590 206360 54640
rect 206140 54520 206150 54590
rect 206350 54520 206360 54590
rect 206140 54480 206360 54520
rect 206140 54410 206150 54480
rect 206350 54410 206360 54480
rect 206140 54360 206360 54410
rect 206640 54590 206860 54640
rect 206640 54520 206650 54590
rect 206850 54520 206860 54590
rect 206640 54480 206860 54520
rect 206640 54410 206650 54480
rect 206850 54410 206860 54480
rect 206640 54360 206860 54410
rect 207140 54590 207360 54640
rect 207140 54520 207150 54590
rect 207350 54520 207360 54590
rect 207140 54480 207360 54520
rect 207140 54410 207150 54480
rect 207350 54410 207360 54480
rect 207140 54360 207360 54410
rect 207640 54590 207860 54640
rect 207640 54520 207650 54590
rect 207850 54520 207860 54590
rect 207640 54480 207860 54520
rect 207640 54410 207650 54480
rect 207850 54410 207860 54480
rect 207640 54360 207860 54410
rect 204000 54350 208000 54360
rect 204000 54150 204020 54350
rect 204090 54150 204410 54350
rect 204480 54150 204520 54350
rect 204590 54150 204910 54350
rect 204980 54150 205020 54350
rect 205090 54150 205410 54350
rect 205480 54150 205520 54350
rect 205590 54150 205910 54350
rect 205980 54150 206020 54350
rect 206090 54150 206410 54350
rect 206480 54150 206520 54350
rect 206590 54150 206910 54350
rect 206980 54150 207020 54350
rect 207090 54150 207410 54350
rect 207480 54150 207520 54350
rect 207590 54150 207910 54350
rect 207980 54150 208000 54350
rect 204000 54140 208000 54150
rect 204140 54090 204360 54140
rect 204140 54020 204150 54090
rect 204350 54020 204360 54090
rect 204140 53980 204360 54020
rect 204140 53910 204150 53980
rect 204350 53910 204360 53980
rect 204140 53860 204360 53910
rect 204640 54090 204860 54140
rect 204640 54020 204650 54090
rect 204850 54020 204860 54090
rect 204640 53980 204860 54020
rect 204640 53910 204650 53980
rect 204850 53910 204860 53980
rect 204640 53860 204860 53910
rect 205140 54090 205360 54140
rect 205140 54020 205150 54090
rect 205350 54020 205360 54090
rect 205140 53980 205360 54020
rect 205140 53910 205150 53980
rect 205350 53910 205360 53980
rect 205140 53860 205360 53910
rect 205640 54090 205860 54140
rect 205640 54020 205650 54090
rect 205850 54020 205860 54090
rect 205640 53980 205860 54020
rect 205640 53910 205650 53980
rect 205850 53910 205860 53980
rect 205640 53860 205860 53910
rect 206140 54090 206360 54140
rect 206140 54020 206150 54090
rect 206350 54020 206360 54090
rect 206140 53980 206360 54020
rect 206140 53910 206150 53980
rect 206350 53910 206360 53980
rect 206140 53860 206360 53910
rect 206640 54090 206860 54140
rect 206640 54020 206650 54090
rect 206850 54020 206860 54090
rect 206640 53980 206860 54020
rect 206640 53910 206650 53980
rect 206850 53910 206860 53980
rect 206640 53860 206860 53910
rect 207140 54090 207360 54140
rect 207140 54020 207150 54090
rect 207350 54020 207360 54090
rect 207140 53980 207360 54020
rect 207140 53910 207150 53980
rect 207350 53910 207360 53980
rect 207140 53860 207360 53910
rect 207640 54090 207860 54140
rect 207640 54020 207650 54090
rect 207850 54020 207860 54090
rect 207640 53980 207860 54020
rect 207640 53910 207650 53980
rect 207850 53910 207860 53980
rect 207640 53860 207860 53910
rect 204000 53850 208000 53860
rect 204000 53650 204020 53850
rect 204090 53650 204410 53850
rect 204480 53650 204520 53850
rect 204590 53650 204910 53850
rect 204980 53650 205020 53850
rect 205090 53650 205410 53850
rect 205480 53650 205520 53850
rect 205590 53650 205910 53850
rect 205980 53650 206020 53850
rect 206090 53650 206410 53850
rect 206480 53650 206520 53850
rect 206590 53650 206910 53850
rect 206980 53650 207020 53850
rect 207090 53650 207410 53850
rect 207480 53650 207520 53850
rect 207590 53650 207910 53850
rect 207980 53650 208000 53850
rect 204000 53640 208000 53650
rect 204140 53590 204360 53640
rect 204140 53520 204150 53590
rect 204350 53520 204360 53590
rect 204140 53480 204360 53520
rect 204140 53410 204150 53480
rect 204350 53410 204360 53480
rect 204140 53360 204360 53410
rect 204640 53590 204860 53640
rect 204640 53520 204650 53590
rect 204850 53520 204860 53590
rect 204640 53480 204860 53520
rect 204640 53410 204650 53480
rect 204850 53410 204860 53480
rect 204640 53360 204860 53410
rect 205140 53590 205360 53640
rect 205140 53520 205150 53590
rect 205350 53520 205360 53590
rect 205140 53480 205360 53520
rect 205140 53410 205150 53480
rect 205350 53410 205360 53480
rect 205140 53360 205360 53410
rect 205640 53590 205860 53640
rect 205640 53520 205650 53590
rect 205850 53520 205860 53590
rect 205640 53480 205860 53520
rect 205640 53410 205650 53480
rect 205850 53410 205860 53480
rect 205640 53360 205860 53410
rect 206140 53590 206360 53640
rect 206140 53520 206150 53590
rect 206350 53520 206360 53590
rect 206140 53480 206360 53520
rect 206140 53410 206150 53480
rect 206350 53410 206360 53480
rect 206140 53360 206360 53410
rect 206640 53590 206860 53640
rect 206640 53520 206650 53590
rect 206850 53520 206860 53590
rect 206640 53480 206860 53520
rect 206640 53410 206650 53480
rect 206850 53410 206860 53480
rect 206640 53360 206860 53410
rect 207140 53590 207360 53640
rect 207140 53520 207150 53590
rect 207350 53520 207360 53590
rect 207140 53480 207360 53520
rect 207140 53410 207150 53480
rect 207350 53410 207360 53480
rect 207140 53360 207360 53410
rect 207640 53590 207860 53640
rect 207640 53520 207650 53590
rect 207850 53520 207860 53590
rect 207640 53480 207860 53520
rect 207640 53410 207650 53480
rect 207850 53410 207860 53480
rect 207640 53360 207860 53410
rect 204000 53350 208000 53360
rect 204000 53150 204020 53350
rect 204090 53150 204410 53350
rect 204480 53150 204520 53350
rect 204590 53150 204910 53350
rect 204980 53150 205020 53350
rect 205090 53150 205410 53350
rect 205480 53150 205520 53350
rect 205590 53150 205910 53350
rect 205980 53150 206020 53350
rect 206090 53150 206410 53350
rect 206480 53150 206520 53350
rect 206590 53150 206910 53350
rect 206980 53150 207020 53350
rect 207090 53150 207410 53350
rect 207480 53150 207520 53350
rect 207590 53150 207910 53350
rect 207980 53150 208000 53350
rect 204000 53140 208000 53150
rect 204140 53090 204360 53140
rect 204140 53020 204150 53090
rect 204350 53020 204360 53090
rect 204140 52980 204360 53020
rect 204140 52910 204150 52980
rect 204350 52910 204360 52980
rect 204140 52860 204360 52910
rect 204640 53090 204860 53140
rect 204640 53020 204650 53090
rect 204850 53020 204860 53090
rect 204640 52980 204860 53020
rect 204640 52910 204650 52980
rect 204850 52910 204860 52980
rect 204640 52860 204860 52910
rect 205140 53090 205360 53140
rect 205140 53020 205150 53090
rect 205350 53020 205360 53090
rect 205140 52980 205360 53020
rect 205140 52910 205150 52980
rect 205350 52910 205360 52980
rect 205140 52860 205360 52910
rect 205640 53090 205860 53140
rect 205640 53020 205650 53090
rect 205850 53020 205860 53090
rect 205640 52980 205860 53020
rect 205640 52910 205650 52980
rect 205850 52910 205860 52980
rect 205640 52860 205860 52910
rect 206140 53090 206360 53140
rect 206140 53020 206150 53090
rect 206350 53020 206360 53090
rect 206140 52980 206360 53020
rect 206140 52910 206150 52980
rect 206350 52910 206360 52980
rect 206140 52860 206360 52910
rect 206640 53090 206860 53140
rect 206640 53020 206650 53090
rect 206850 53020 206860 53090
rect 206640 52980 206860 53020
rect 206640 52910 206650 52980
rect 206850 52910 206860 52980
rect 206640 52860 206860 52910
rect 207140 53090 207360 53140
rect 207140 53020 207150 53090
rect 207350 53020 207360 53090
rect 207140 52980 207360 53020
rect 207140 52910 207150 52980
rect 207350 52910 207360 52980
rect 207140 52860 207360 52910
rect 207640 53090 207860 53140
rect 207640 53020 207650 53090
rect 207850 53020 207860 53090
rect 207640 52980 207860 53020
rect 207640 52910 207650 52980
rect 207850 52910 207860 52980
rect 207640 52860 207860 52910
rect 204000 52850 208000 52860
rect 204000 52650 204020 52850
rect 204090 52650 204410 52850
rect 204480 52650 204520 52850
rect 204590 52650 204910 52850
rect 204980 52650 205020 52850
rect 205090 52650 205410 52850
rect 205480 52650 205520 52850
rect 205590 52650 205910 52850
rect 205980 52650 206020 52850
rect 206090 52650 206410 52850
rect 206480 52650 206520 52850
rect 206590 52650 206910 52850
rect 206980 52650 207020 52850
rect 207090 52650 207410 52850
rect 207480 52650 207520 52850
rect 207590 52650 207910 52850
rect 207980 52650 208000 52850
rect 204000 52640 208000 52650
rect 204140 52590 204360 52640
rect 204140 52520 204150 52590
rect 204350 52520 204360 52590
rect 204140 52480 204360 52520
rect 204140 52410 204150 52480
rect 204350 52410 204360 52480
rect 204140 52360 204360 52410
rect 204640 52590 204860 52640
rect 204640 52520 204650 52590
rect 204850 52520 204860 52590
rect 204640 52480 204860 52520
rect 204640 52410 204650 52480
rect 204850 52410 204860 52480
rect 204640 52360 204860 52410
rect 205140 52590 205360 52640
rect 205140 52520 205150 52590
rect 205350 52520 205360 52590
rect 205140 52480 205360 52520
rect 205140 52410 205150 52480
rect 205350 52410 205360 52480
rect 205140 52360 205360 52410
rect 205640 52590 205860 52640
rect 205640 52520 205650 52590
rect 205850 52520 205860 52590
rect 205640 52480 205860 52520
rect 205640 52410 205650 52480
rect 205850 52410 205860 52480
rect 205640 52360 205860 52410
rect 206140 52590 206360 52640
rect 206140 52520 206150 52590
rect 206350 52520 206360 52590
rect 206140 52480 206360 52520
rect 206140 52410 206150 52480
rect 206350 52410 206360 52480
rect 206140 52360 206360 52410
rect 206640 52590 206860 52640
rect 206640 52520 206650 52590
rect 206850 52520 206860 52590
rect 206640 52480 206860 52520
rect 206640 52410 206650 52480
rect 206850 52410 206860 52480
rect 206640 52360 206860 52410
rect 207140 52590 207360 52640
rect 207140 52520 207150 52590
rect 207350 52520 207360 52590
rect 207140 52480 207360 52520
rect 207140 52410 207150 52480
rect 207350 52410 207360 52480
rect 207140 52360 207360 52410
rect 207640 52590 207860 52640
rect 207640 52520 207650 52590
rect 207850 52520 207860 52590
rect 207640 52480 207860 52520
rect 207640 52410 207650 52480
rect 207850 52410 207860 52480
rect 207640 52360 207860 52410
rect 204000 52350 208000 52360
rect 204000 52150 204020 52350
rect 204090 52150 204410 52350
rect 204480 52150 204520 52350
rect 204590 52150 204910 52350
rect 204980 52150 205020 52350
rect 205090 52150 205410 52350
rect 205480 52150 205520 52350
rect 205590 52150 205910 52350
rect 205980 52150 206020 52350
rect 206090 52150 206410 52350
rect 206480 52150 206520 52350
rect 206590 52150 206910 52350
rect 206980 52150 207020 52350
rect 207090 52150 207410 52350
rect 207480 52150 207520 52350
rect 207590 52150 207910 52350
rect 207980 52150 208000 52350
rect 204000 52140 208000 52150
rect 204140 52090 204360 52140
rect 204140 52020 204150 52090
rect 204350 52020 204360 52090
rect 204140 51980 204360 52020
rect 204140 51910 204150 51980
rect 204350 51910 204360 51980
rect 204140 51860 204360 51910
rect 204640 52090 204860 52140
rect 204640 52020 204650 52090
rect 204850 52020 204860 52090
rect 204640 51980 204860 52020
rect 204640 51910 204650 51980
rect 204850 51910 204860 51980
rect 204640 51860 204860 51910
rect 205140 52090 205360 52140
rect 205140 52020 205150 52090
rect 205350 52020 205360 52090
rect 205140 51980 205360 52020
rect 205140 51910 205150 51980
rect 205350 51910 205360 51980
rect 205140 51860 205360 51910
rect 205640 52090 205860 52140
rect 205640 52020 205650 52090
rect 205850 52020 205860 52090
rect 205640 51980 205860 52020
rect 205640 51910 205650 51980
rect 205850 51910 205860 51980
rect 205640 51860 205860 51910
rect 206140 52090 206360 52140
rect 206140 52020 206150 52090
rect 206350 52020 206360 52090
rect 206140 51980 206360 52020
rect 206140 51910 206150 51980
rect 206350 51910 206360 51980
rect 206140 51860 206360 51910
rect 206640 52090 206860 52140
rect 206640 52020 206650 52090
rect 206850 52020 206860 52090
rect 206640 51980 206860 52020
rect 206640 51910 206650 51980
rect 206850 51910 206860 51980
rect 206640 51860 206860 51910
rect 207140 52090 207360 52140
rect 207140 52020 207150 52090
rect 207350 52020 207360 52090
rect 207140 51980 207360 52020
rect 207140 51910 207150 51980
rect 207350 51910 207360 51980
rect 207140 51860 207360 51910
rect 207640 52090 207860 52140
rect 207640 52020 207650 52090
rect 207850 52020 207860 52090
rect 207640 51980 207860 52020
rect 207640 51910 207650 51980
rect 207850 51910 207860 51980
rect 207640 51860 207860 51910
rect 204000 51850 208000 51860
rect 204000 51650 204020 51850
rect 204090 51650 204410 51850
rect 204480 51650 204520 51850
rect 204590 51650 204910 51850
rect 204980 51650 205020 51850
rect 205090 51650 205410 51850
rect 205480 51650 205520 51850
rect 205590 51650 205910 51850
rect 205980 51650 206020 51850
rect 206090 51650 206410 51850
rect 206480 51650 206520 51850
rect 206590 51650 206910 51850
rect 206980 51650 207020 51850
rect 207090 51650 207410 51850
rect 207480 51650 207520 51850
rect 207590 51650 207910 51850
rect 207980 51650 208000 51850
rect 204000 51640 208000 51650
rect 204140 51590 204360 51640
rect 204140 51520 204150 51590
rect 204350 51520 204360 51590
rect 204140 51480 204360 51520
rect 204140 51410 204150 51480
rect 204350 51410 204360 51480
rect 204140 51360 204360 51410
rect 204640 51590 204860 51640
rect 204640 51520 204650 51590
rect 204850 51520 204860 51590
rect 204640 51480 204860 51520
rect 204640 51410 204650 51480
rect 204850 51410 204860 51480
rect 204640 51360 204860 51410
rect 205140 51590 205360 51640
rect 205140 51520 205150 51590
rect 205350 51520 205360 51590
rect 205140 51480 205360 51520
rect 205140 51410 205150 51480
rect 205350 51410 205360 51480
rect 205140 51360 205360 51410
rect 205640 51590 205860 51640
rect 205640 51520 205650 51590
rect 205850 51520 205860 51590
rect 205640 51480 205860 51520
rect 205640 51410 205650 51480
rect 205850 51410 205860 51480
rect 205640 51360 205860 51410
rect 206140 51590 206360 51640
rect 206140 51520 206150 51590
rect 206350 51520 206360 51590
rect 206140 51480 206360 51520
rect 206140 51410 206150 51480
rect 206350 51410 206360 51480
rect 206140 51360 206360 51410
rect 206640 51590 206860 51640
rect 206640 51520 206650 51590
rect 206850 51520 206860 51590
rect 206640 51480 206860 51520
rect 206640 51410 206650 51480
rect 206850 51410 206860 51480
rect 206640 51360 206860 51410
rect 207140 51590 207360 51640
rect 207140 51520 207150 51590
rect 207350 51520 207360 51590
rect 207140 51480 207360 51520
rect 207140 51410 207150 51480
rect 207350 51410 207360 51480
rect 207140 51360 207360 51410
rect 207640 51590 207860 51640
rect 207640 51520 207650 51590
rect 207850 51520 207860 51590
rect 207640 51480 207860 51520
rect 207640 51410 207650 51480
rect 207850 51410 207860 51480
rect 207640 51360 207860 51410
rect 204000 51350 208000 51360
rect 204000 51150 204020 51350
rect 204090 51150 204410 51350
rect 204480 51150 204520 51350
rect 204590 51150 204910 51350
rect 204980 51150 205020 51350
rect 205090 51150 205410 51350
rect 205480 51150 205520 51350
rect 205590 51150 205910 51350
rect 205980 51150 206020 51350
rect 206090 51150 206410 51350
rect 206480 51150 206520 51350
rect 206590 51150 206910 51350
rect 206980 51150 207020 51350
rect 207090 51150 207410 51350
rect 207480 51150 207520 51350
rect 207590 51150 207910 51350
rect 207980 51150 208000 51350
rect 204000 51140 208000 51150
rect 204140 51090 204360 51140
rect 204140 51020 204150 51090
rect 204350 51020 204360 51090
rect 204140 50980 204360 51020
rect 204140 50910 204150 50980
rect 204350 50910 204360 50980
rect 204140 50860 204360 50910
rect 204640 51090 204860 51140
rect 204640 51020 204650 51090
rect 204850 51020 204860 51090
rect 204640 50980 204860 51020
rect 204640 50910 204650 50980
rect 204850 50910 204860 50980
rect 204640 50860 204860 50910
rect 205140 51090 205360 51140
rect 205140 51020 205150 51090
rect 205350 51020 205360 51090
rect 205140 50980 205360 51020
rect 205140 50910 205150 50980
rect 205350 50910 205360 50980
rect 205140 50860 205360 50910
rect 205640 51090 205860 51140
rect 205640 51020 205650 51090
rect 205850 51020 205860 51090
rect 205640 50980 205860 51020
rect 205640 50910 205650 50980
rect 205850 50910 205860 50980
rect 205640 50860 205860 50910
rect 206140 51090 206360 51140
rect 206140 51020 206150 51090
rect 206350 51020 206360 51090
rect 206140 50980 206360 51020
rect 206140 50910 206150 50980
rect 206350 50910 206360 50980
rect 206140 50860 206360 50910
rect 206640 51090 206860 51140
rect 206640 51020 206650 51090
rect 206850 51020 206860 51090
rect 206640 50980 206860 51020
rect 206640 50910 206650 50980
rect 206850 50910 206860 50980
rect 206640 50860 206860 50910
rect 207140 51090 207360 51140
rect 207140 51020 207150 51090
rect 207350 51020 207360 51090
rect 207140 50980 207360 51020
rect 207140 50910 207150 50980
rect 207350 50910 207360 50980
rect 207140 50860 207360 50910
rect 207640 51090 207860 51140
rect 207640 51020 207650 51090
rect 207850 51020 207860 51090
rect 207640 50980 207860 51020
rect 207640 50910 207650 50980
rect 207850 50910 207860 50980
rect 207640 50860 207860 50910
rect 204000 50850 208000 50860
rect 204000 50650 204020 50850
rect 204090 50650 204410 50850
rect 204480 50650 204520 50850
rect 204590 50650 204910 50850
rect 204980 50650 205020 50850
rect 205090 50650 205410 50850
rect 205480 50650 205520 50850
rect 205590 50650 205910 50850
rect 205980 50650 206020 50850
rect 206090 50650 206410 50850
rect 206480 50650 206520 50850
rect 206590 50650 206910 50850
rect 206980 50650 207020 50850
rect 207090 50650 207410 50850
rect 207480 50650 207520 50850
rect 207590 50650 207910 50850
rect 207980 50650 208000 50850
rect 204000 50640 208000 50650
rect 204140 50590 204360 50640
rect 204140 50520 204150 50590
rect 204350 50520 204360 50590
rect 204140 50480 204360 50520
rect 204140 50410 204150 50480
rect 204350 50410 204360 50480
rect 204140 50360 204360 50410
rect 204640 50590 204860 50640
rect 204640 50520 204650 50590
rect 204850 50520 204860 50590
rect 204640 50480 204860 50520
rect 204640 50410 204650 50480
rect 204850 50410 204860 50480
rect 204640 50360 204860 50410
rect 205140 50590 205360 50640
rect 205140 50520 205150 50590
rect 205350 50520 205360 50590
rect 205140 50480 205360 50520
rect 205140 50410 205150 50480
rect 205350 50410 205360 50480
rect 205140 50360 205360 50410
rect 205640 50590 205860 50640
rect 205640 50520 205650 50590
rect 205850 50520 205860 50590
rect 205640 50480 205860 50520
rect 205640 50410 205650 50480
rect 205850 50410 205860 50480
rect 205640 50360 205860 50410
rect 206140 50590 206360 50640
rect 206140 50520 206150 50590
rect 206350 50520 206360 50590
rect 206140 50480 206360 50520
rect 206140 50410 206150 50480
rect 206350 50410 206360 50480
rect 206140 50360 206360 50410
rect 206640 50590 206860 50640
rect 206640 50520 206650 50590
rect 206850 50520 206860 50590
rect 206640 50480 206860 50520
rect 206640 50410 206650 50480
rect 206850 50410 206860 50480
rect 206640 50360 206860 50410
rect 207140 50590 207360 50640
rect 207140 50520 207150 50590
rect 207350 50520 207360 50590
rect 207140 50480 207360 50520
rect 207140 50410 207150 50480
rect 207350 50410 207360 50480
rect 207140 50360 207360 50410
rect 207640 50590 207860 50640
rect 207640 50520 207650 50590
rect 207850 50520 207860 50590
rect 207640 50480 207860 50520
rect 207640 50410 207650 50480
rect 207850 50410 207860 50480
rect 207640 50360 207860 50410
rect 204000 50350 208000 50360
rect 204000 50150 204020 50350
rect 204090 50150 204410 50350
rect 204480 50150 204520 50350
rect 204590 50150 204910 50350
rect 204980 50150 205020 50350
rect 205090 50150 205410 50350
rect 205480 50150 205520 50350
rect 205590 50150 205910 50350
rect 205980 50150 206020 50350
rect 206090 50150 206410 50350
rect 206480 50150 206520 50350
rect 206590 50150 206910 50350
rect 206980 50150 207020 50350
rect 207090 50150 207410 50350
rect 207480 50150 207520 50350
rect 207590 50150 207910 50350
rect 207980 50150 208000 50350
rect 204000 50140 208000 50150
rect 204140 50090 204360 50140
rect 204140 50020 204150 50090
rect 204350 50020 204360 50090
rect 204140 49980 204360 50020
rect 204140 49910 204150 49980
rect 204350 49910 204360 49980
rect 204140 49860 204360 49910
rect 204640 50090 204860 50140
rect 204640 50020 204650 50090
rect 204850 50020 204860 50090
rect 204640 49980 204860 50020
rect 204640 49910 204650 49980
rect 204850 49910 204860 49980
rect 204640 49860 204860 49910
rect 205140 50090 205360 50140
rect 205140 50020 205150 50090
rect 205350 50020 205360 50090
rect 205140 49980 205360 50020
rect 205140 49910 205150 49980
rect 205350 49910 205360 49980
rect 205140 49860 205360 49910
rect 205640 50090 205860 50140
rect 205640 50020 205650 50090
rect 205850 50020 205860 50090
rect 205640 49980 205860 50020
rect 205640 49910 205650 49980
rect 205850 49910 205860 49980
rect 205640 49860 205860 49910
rect 206140 50090 206360 50140
rect 206140 50020 206150 50090
rect 206350 50020 206360 50090
rect 206140 49980 206360 50020
rect 206140 49910 206150 49980
rect 206350 49910 206360 49980
rect 206140 49860 206360 49910
rect 206640 50090 206860 50140
rect 206640 50020 206650 50090
rect 206850 50020 206860 50090
rect 206640 49980 206860 50020
rect 206640 49910 206650 49980
rect 206850 49910 206860 49980
rect 206640 49860 206860 49910
rect 207140 50090 207360 50140
rect 207140 50020 207150 50090
rect 207350 50020 207360 50090
rect 207140 49980 207360 50020
rect 207140 49910 207150 49980
rect 207350 49910 207360 49980
rect 207140 49860 207360 49910
rect 207640 50090 207860 50140
rect 207640 50020 207650 50090
rect 207850 50020 207860 50090
rect 207640 49980 207860 50020
rect 207640 49910 207650 49980
rect 207850 49910 207860 49980
rect 207640 49860 207860 49910
rect 204000 49850 208000 49860
rect 204000 49650 204020 49850
rect 204090 49650 204410 49850
rect 204480 49650 204520 49850
rect 204590 49650 204910 49850
rect 204980 49650 205020 49850
rect 205090 49650 205410 49850
rect 205480 49650 205520 49850
rect 205590 49650 205910 49850
rect 205980 49650 206020 49850
rect 206090 49650 206410 49850
rect 206480 49650 206520 49850
rect 206590 49650 206910 49850
rect 206980 49650 207020 49850
rect 207090 49650 207410 49850
rect 207480 49650 207520 49850
rect 207590 49650 207910 49850
rect 207980 49650 208000 49850
rect 204000 49640 208000 49650
rect 204140 49590 204360 49640
rect 204140 49520 204150 49590
rect 204350 49520 204360 49590
rect 204140 49480 204360 49520
rect 204140 49410 204150 49480
rect 204350 49410 204360 49480
rect 204140 49360 204360 49410
rect 204640 49590 204860 49640
rect 204640 49520 204650 49590
rect 204850 49520 204860 49590
rect 204640 49480 204860 49520
rect 204640 49410 204650 49480
rect 204850 49410 204860 49480
rect 204640 49360 204860 49410
rect 205140 49590 205360 49640
rect 205140 49520 205150 49590
rect 205350 49520 205360 49590
rect 205140 49480 205360 49520
rect 205140 49410 205150 49480
rect 205350 49410 205360 49480
rect 205140 49360 205360 49410
rect 205640 49590 205860 49640
rect 205640 49520 205650 49590
rect 205850 49520 205860 49590
rect 205640 49480 205860 49520
rect 205640 49410 205650 49480
rect 205850 49410 205860 49480
rect 205640 49360 205860 49410
rect 206140 49590 206360 49640
rect 206140 49520 206150 49590
rect 206350 49520 206360 49590
rect 206140 49480 206360 49520
rect 206140 49410 206150 49480
rect 206350 49410 206360 49480
rect 206140 49360 206360 49410
rect 206640 49590 206860 49640
rect 206640 49520 206650 49590
rect 206850 49520 206860 49590
rect 206640 49480 206860 49520
rect 206640 49410 206650 49480
rect 206850 49410 206860 49480
rect 206640 49360 206860 49410
rect 207140 49590 207360 49640
rect 207140 49520 207150 49590
rect 207350 49520 207360 49590
rect 207140 49480 207360 49520
rect 207140 49410 207150 49480
rect 207350 49410 207360 49480
rect 207140 49360 207360 49410
rect 207640 49590 207860 49640
rect 207640 49520 207650 49590
rect 207850 49520 207860 49590
rect 207640 49480 207860 49520
rect 207640 49410 207650 49480
rect 207850 49410 207860 49480
rect 207640 49360 207860 49410
rect 204000 49350 208000 49360
rect 204000 49150 204020 49350
rect 204090 49150 204410 49350
rect 204480 49150 204520 49350
rect 204590 49150 204910 49350
rect 204980 49150 205020 49350
rect 205090 49150 205410 49350
rect 205480 49150 205520 49350
rect 205590 49150 205910 49350
rect 205980 49150 206020 49350
rect 206090 49150 206410 49350
rect 206480 49150 206520 49350
rect 206590 49150 206910 49350
rect 206980 49150 207020 49350
rect 207090 49150 207410 49350
rect 207480 49150 207520 49350
rect 207590 49150 207910 49350
rect 207980 49150 208000 49350
rect 204000 49140 208000 49150
rect 204140 49090 204360 49140
rect 204140 49020 204150 49090
rect 204350 49020 204360 49090
rect 204140 48980 204360 49020
rect 204140 48910 204150 48980
rect 204350 48910 204360 48980
rect 204140 48860 204360 48910
rect 204640 49090 204860 49140
rect 204640 49020 204650 49090
rect 204850 49020 204860 49090
rect 204640 48980 204860 49020
rect 204640 48910 204650 48980
rect 204850 48910 204860 48980
rect 204640 48860 204860 48910
rect 205140 49090 205360 49140
rect 205140 49020 205150 49090
rect 205350 49020 205360 49090
rect 205140 48980 205360 49020
rect 205140 48910 205150 48980
rect 205350 48910 205360 48980
rect 205140 48860 205360 48910
rect 205640 49090 205860 49140
rect 205640 49020 205650 49090
rect 205850 49020 205860 49090
rect 205640 48980 205860 49020
rect 205640 48910 205650 48980
rect 205850 48910 205860 48980
rect 205640 48860 205860 48910
rect 206140 49090 206360 49140
rect 206140 49020 206150 49090
rect 206350 49020 206360 49090
rect 206140 48980 206360 49020
rect 206140 48910 206150 48980
rect 206350 48910 206360 48980
rect 206140 48860 206360 48910
rect 206640 49090 206860 49140
rect 206640 49020 206650 49090
rect 206850 49020 206860 49090
rect 206640 48980 206860 49020
rect 206640 48910 206650 48980
rect 206850 48910 206860 48980
rect 206640 48860 206860 48910
rect 207140 49090 207360 49140
rect 207140 49020 207150 49090
rect 207350 49020 207360 49090
rect 207140 48980 207360 49020
rect 207140 48910 207150 48980
rect 207350 48910 207360 48980
rect 207140 48860 207360 48910
rect 207640 49090 207860 49140
rect 207640 49020 207650 49090
rect 207850 49020 207860 49090
rect 207640 48980 207860 49020
rect 207640 48910 207650 48980
rect 207850 48910 207860 48980
rect 207640 48860 207860 48910
rect 204000 48850 208000 48860
rect 204000 48650 204020 48850
rect 204090 48650 204410 48850
rect 204480 48650 204520 48850
rect 204590 48650 204910 48850
rect 204980 48650 205020 48850
rect 205090 48650 205410 48850
rect 205480 48650 205520 48850
rect 205590 48650 205910 48850
rect 205980 48650 206020 48850
rect 206090 48650 206410 48850
rect 206480 48650 206520 48850
rect 206590 48650 206910 48850
rect 206980 48650 207020 48850
rect 207090 48650 207410 48850
rect 207480 48650 207520 48850
rect 207590 48650 207910 48850
rect 207980 48650 208000 48850
rect 204000 48640 208000 48650
rect 204140 48590 204360 48640
rect 204140 48520 204150 48590
rect 204350 48520 204360 48590
rect 204140 48480 204360 48520
rect 204140 48410 204150 48480
rect 204350 48410 204360 48480
rect 204140 48360 204360 48410
rect 204640 48590 204860 48640
rect 204640 48520 204650 48590
rect 204850 48520 204860 48590
rect 204640 48480 204860 48520
rect 204640 48410 204650 48480
rect 204850 48410 204860 48480
rect 204640 48360 204860 48410
rect 205140 48590 205360 48640
rect 205140 48520 205150 48590
rect 205350 48520 205360 48590
rect 205140 48480 205360 48520
rect 205140 48410 205150 48480
rect 205350 48410 205360 48480
rect 205140 48360 205360 48410
rect 205640 48590 205860 48640
rect 205640 48520 205650 48590
rect 205850 48520 205860 48590
rect 205640 48480 205860 48520
rect 205640 48410 205650 48480
rect 205850 48410 205860 48480
rect 205640 48360 205860 48410
rect 206140 48590 206360 48640
rect 206140 48520 206150 48590
rect 206350 48520 206360 48590
rect 206140 48480 206360 48520
rect 206140 48410 206150 48480
rect 206350 48410 206360 48480
rect 206140 48360 206360 48410
rect 206640 48590 206860 48640
rect 206640 48520 206650 48590
rect 206850 48520 206860 48590
rect 206640 48480 206860 48520
rect 206640 48410 206650 48480
rect 206850 48410 206860 48480
rect 206640 48360 206860 48410
rect 207140 48590 207360 48640
rect 207140 48520 207150 48590
rect 207350 48520 207360 48590
rect 207140 48480 207360 48520
rect 207140 48410 207150 48480
rect 207350 48410 207360 48480
rect 207140 48360 207360 48410
rect 207640 48590 207860 48640
rect 207640 48520 207650 48590
rect 207850 48520 207860 48590
rect 207640 48480 207860 48520
rect 207640 48410 207650 48480
rect 207850 48410 207860 48480
rect 207640 48360 207860 48410
rect 204000 48350 208000 48360
rect 204000 48150 204020 48350
rect 204090 48150 204410 48350
rect 204480 48150 204520 48350
rect 204590 48150 204910 48350
rect 204980 48150 205020 48350
rect 205090 48150 205410 48350
rect 205480 48150 205520 48350
rect 205590 48150 205910 48350
rect 205980 48150 206020 48350
rect 206090 48150 206410 48350
rect 206480 48150 206520 48350
rect 206590 48150 206910 48350
rect 206980 48150 207020 48350
rect 207090 48150 207410 48350
rect 207480 48150 207520 48350
rect 207590 48150 207910 48350
rect 207980 48150 208000 48350
rect 204000 48140 208000 48150
rect 204140 48090 204360 48140
rect 204140 48020 204150 48090
rect 204350 48020 204360 48090
rect 204140 47980 204360 48020
rect 204140 47910 204150 47980
rect 204350 47910 204360 47980
rect 204140 47860 204360 47910
rect 204640 48090 204860 48140
rect 204640 48020 204650 48090
rect 204850 48020 204860 48090
rect 204640 47980 204860 48020
rect 204640 47910 204650 47980
rect 204850 47910 204860 47980
rect 204640 47860 204860 47910
rect 205140 48090 205360 48140
rect 205140 48020 205150 48090
rect 205350 48020 205360 48090
rect 205140 47980 205360 48020
rect 205140 47910 205150 47980
rect 205350 47910 205360 47980
rect 205140 47860 205360 47910
rect 205640 48090 205860 48140
rect 205640 48020 205650 48090
rect 205850 48020 205860 48090
rect 205640 47980 205860 48020
rect 205640 47910 205650 47980
rect 205850 47910 205860 47980
rect 205640 47860 205860 47910
rect 206140 48090 206360 48140
rect 206140 48020 206150 48090
rect 206350 48020 206360 48090
rect 206140 47980 206360 48020
rect 206140 47910 206150 47980
rect 206350 47910 206360 47980
rect 206140 47860 206360 47910
rect 206640 48090 206860 48140
rect 206640 48020 206650 48090
rect 206850 48020 206860 48090
rect 206640 47980 206860 48020
rect 206640 47910 206650 47980
rect 206850 47910 206860 47980
rect 206640 47860 206860 47910
rect 207140 48090 207360 48140
rect 207140 48020 207150 48090
rect 207350 48020 207360 48090
rect 207140 47980 207360 48020
rect 207140 47910 207150 47980
rect 207350 47910 207360 47980
rect 207140 47860 207360 47910
rect 207640 48090 207860 48140
rect 207640 48020 207650 48090
rect 207850 48020 207860 48090
rect 207640 47980 207860 48020
rect 207640 47910 207650 47980
rect 207850 47910 207860 47980
rect 207640 47860 207860 47910
rect 204000 47850 208000 47860
rect 204000 47650 204020 47850
rect 204090 47650 204410 47850
rect 204480 47650 204520 47850
rect 204590 47650 204910 47850
rect 204980 47650 205020 47850
rect 205090 47650 205410 47850
rect 205480 47650 205520 47850
rect 205590 47650 205910 47850
rect 205980 47650 206020 47850
rect 206090 47650 206410 47850
rect 206480 47650 206520 47850
rect 206590 47650 206910 47850
rect 206980 47650 207020 47850
rect 207090 47650 207410 47850
rect 207480 47650 207520 47850
rect 207590 47650 207910 47850
rect 207980 47650 208000 47850
rect 204000 47640 208000 47650
rect 204140 47590 204360 47640
rect 204140 47520 204150 47590
rect 204350 47520 204360 47590
rect 204140 47480 204360 47520
rect 204140 47410 204150 47480
rect 204350 47410 204360 47480
rect 204140 47360 204360 47410
rect 204640 47590 204860 47640
rect 204640 47520 204650 47590
rect 204850 47520 204860 47590
rect 204640 47480 204860 47520
rect 204640 47410 204650 47480
rect 204850 47410 204860 47480
rect 204640 47360 204860 47410
rect 205140 47590 205360 47640
rect 205140 47520 205150 47590
rect 205350 47520 205360 47590
rect 205140 47480 205360 47520
rect 205140 47410 205150 47480
rect 205350 47410 205360 47480
rect 205140 47360 205360 47410
rect 205640 47590 205860 47640
rect 205640 47520 205650 47590
rect 205850 47520 205860 47590
rect 205640 47480 205860 47520
rect 205640 47410 205650 47480
rect 205850 47410 205860 47480
rect 205640 47360 205860 47410
rect 206140 47590 206360 47640
rect 206140 47520 206150 47590
rect 206350 47520 206360 47590
rect 206140 47480 206360 47520
rect 206140 47410 206150 47480
rect 206350 47410 206360 47480
rect 206140 47360 206360 47410
rect 206640 47590 206860 47640
rect 206640 47520 206650 47590
rect 206850 47520 206860 47590
rect 206640 47480 206860 47520
rect 206640 47410 206650 47480
rect 206850 47410 206860 47480
rect 206640 47360 206860 47410
rect 207140 47590 207360 47640
rect 207140 47520 207150 47590
rect 207350 47520 207360 47590
rect 207140 47480 207360 47520
rect 207140 47410 207150 47480
rect 207350 47410 207360 47480
rect 207140 47360 207360 47410
rect 207640 47590 207860 47640
rect 207640 47520 207650 47590
rect 207850 47520 207860 47590
rect 207640 47480 207860 47520
rect 207640 47410 207650 47480
rect 207850 47410 207860 47480
rect 207640 47360 207860 47410
rect 204000 47350 208000 47360
rect 204000 47150 204020 47350
rect 204090 47150 204410 47350
rect 204480 47150 204520 47350
rect 204590 47150 204910 47350
rect 204980 47150 205020 47350
rect 205090 47150 205410 47350
rect 205480 47150 205520 47350
rect 205590 47150 205910 47350
rect 205980 47150 206020 47350
rect 206090 47150 206410 47350
rect 206480 47150 206520 47350
rect 206590 47150 206910 47350
rect 206980 47150 207020 47350
rect 207090 47150 207410 47350
rect 207480 47150 207520 47350
rect 207590 47150 207910 47350
rect 207980 47150 208000 47350
rect 204000 47140 208000 47150
rect 204140 47090 204360 47140
rect 204140 47020 204150 47090
rect 204350 47020 204360 47090
rect 204140 46980 204360 47020
rect 204140 46910 204150 46980
rect 204350 46910 204360 46980
rect 204140 46860 204360 46910
rect 204640 47090 204860 47140
rect 204640 47020 204650 47090
rect 204850 47020 204860 47090
rect 204640 46980 204860 47020
rect 204640 46910 204650 46980
rect 204850 46910 204860 46980
rect 204640 46860 204860 46910
rect 205140 47090 205360 47140
rect 205140 47020 205150 47090
rect 205350 47020 205360 47090
rect 205140 46980 205360 47020
rect 205140 46910 205150 46980
rect 205350 46910 205360 46980
rect 205140 46860 205360 46910
rect 205640 47090 205860 47140
rect 205640 47020 205650 47090
rect 205850 47020 205860 47090
rect 205640 46980 205860 47020
rect 205640 46910 205650 46980
rect 205850 46910 205860 46980
rect 205640 46860 205860 46910
rect 206140 47090 206360 47140
rect 206140 47020 206150 47090
rect 206350 47020 206360 47090
rect 206140 46980 206360 47020
rect 206140 46910 206150 46980
rect 206350 46910 206360 46980
rect 206140 46860 206360 46910
rect 206640 47090 206860 47140
rect 206640 47020 206650 47090
rect 206850 47020 206860 47090
rect 206640 46980 206860 47020
rect 206640 46910 206650 46980
rect 206850 46910 206860 46980
rect 206640 46860 206860 46910
rect 207140 47090 207360 47140
rect 207140 47020 207150 47090
rect 207350 47020 207360 47090
rect 207140 46980 207360 47020
rect 207140 46910 207150 46980
rect 207350 46910 207360 46980
rect 207140 46860 207360 46910
rect 207640 47090 207860 47140
rect 207640 47020 207650 47090
rect 207850 47020 207860 47090
rect 207640 46980 207860 47020
rect 207640 46910 207650 46980
rect 207850 46910 207860 46980
rect 207640 46860 207860 46910
rect 204000 46850 208000 46860
rect 204000 46650 204020 46850
rect 204090 46650 204410 46850
rect 204480 46650 204520 46850
rect 204590 46650 204910 46850
rect 204980 46650 205020 46850
rect 205090 46650 205410 46850
rect 205480 46650 205520 46850
rect 205590 46650 205910 46850
rect 205980 46650 206020 46850
rect 206090 46650 206410 46850
rect 206480 46650 206520 46850
rect 206590 46650 206910 46850
rect 206980 46650 207020 46850
rect 207090 46650 207410 46850
rect 207480 46650 207520 46850
rect 207590 46650 207910 46850
rect 207980 46650 208000 46850
rect 204000 46640 208000 46650
rect 204140 46590 204360 46640
rect 204140 46520 204150 46590
rect 204350 46520 204360 46590
rect 204140 46480 204360 46520
rect 204140 46410 204150 46480
rect 204350 46410 204360 46480
rect 204140 46360 204360 46410
rect 204640 46590 204860 46640
rect 204640 46520 204650 46590
rect 204850 46520 204860 46590
rect 204640 46480 204860 46520
rect 204640 46410 204650 46480
rect 204850 46410 204860 46480
rect 204640 46360 204860 46410
rect 205140 46590 205360 46640
rect 205140 46520 205150 46590
rect 205350 46520 205360 46590
rect 205140 46480 205360 46520
rect 205140 46410 205150 46480
rect 205350 46410 205360 46480
rect 205140 46360 205360 46410
rect 205640 46590 205860 46640
rect 205640 46520 205650 46590
rect 205850 46520 205860 46590
rect 205640 46480 205860 46520
rect 205640 46410 205650 46480
rect 205850 46410 205860 46480
rect 205640 46360 205860 46410
rect 206140 46590 206360 46640
rect 206140 46520 206150 46590
rect 206350 46520 206360 46590
rect 206140 46480 206360 46520
rect 206140 46410 206150 46480
rect 206350 46410 206360 46480
rect 206140 46360 206360 46410
rect 206640 46590 206860 46640
rect 206640 46520 206650 46590
rect 206850 46520 206860 46590
rect 206640 46480 206860 46520
rect 206640 46410 206650 46480
rect 206850 46410 206860 46480
rect 206640 46360 206860 46410
rect 207140 46590 207360 46640
rect 207140 46520 207150 46590
rect 207350 46520 207360 46590
rect 207140 46480 207360 46520
rect 207140 46410 207150 46480
rect 207350 46410 207360 46480
rect 207140 46360 207360 46410
rect 207640 46590 207860 46640
rect 207640 46520 207650 46590
rect 207850 46520 207860 46590
rect 207640 46480 207860 46520
rect 207640 46410 207650 46480
rect 207850 46410 207860 46480
rect 207640 46360 207860 46410
rect 204000 46350 208000 46360
rect 204000 46150 204020 46350
rect 204090 46150 204410 46350
rect 204480 46150 204520 46350
rect 204590 46150 204910 46350
rect 204980 46150 205020 46350
rect 205090 46150 205410 46350
rect 205480 46150 205520 46350
rect 205590 46150 205910 46350
rect 205980 46150 206020 46350
rect 206090 46150 206410 46350
rect 206480 46150 206520 46350
rect 206590 46150 206910 46350
rect 206980 46150 207020 46350
rect 207090 46150 207410 46350
rect 207480 46150 207520 46350
rect 207590 46150 207910 46350
rect 207980 46150 208000 46350
rect 204000 46140 208000 46150
rect 204140 46090 204360 46140
rect 204140 46020 204150 46090
rect 204350 46020 204360 46090
rect 204140 45980 204360 46020
rect 204140 45910 204150 45980
rect 204350 45910 204360 45980
rect 204140 45860 204360 45910
rect 204640 46090 204860 46140
rect 204640 46020 204650 46090
rect 204850 46020 204860 46090
rect 204640 45980 204860 46020
rect 204640 45910 204650 45980
rect 204850 45910 204860 45980
rect 204640 45860 204860 45910
rect 205140 46090 205360 46140
rect 205140 46020 205150 46090
rect 205350 46020 205360 46090
rect 205140 45980 205360 46020
rect 205140 45910 205150 45980
rect 205350 45910 205360 45980
rect 205140 45860 205360 45910
rect 205640 46090 205860 46140
rect 205640 46020 205650 46090
rect 205850 46020 205860 46090
rect 205640 45980 205860 46020
rect 205640 45910 205650 45980
rect 205850 45910 205860 45980
rect 205640 45860 205860 45910
rect 206140 46090 206360 46140
rect 206140 46020 206150 46090
rect 206350 46020 206360 46090
rect 206140 45980 206360 46020
rect 206140 45910 206150 45980
rect 206350 45910 206360 45980
rect 206140 45860 206360 45910
rect 206640 46090 206860 46140
rect 206640 46020 206650 46090
rect 206850 46020 206860 46090
rect 206640 45980 206860 46020
rect 206640 45910 206650 45980
rect 206850 45910 206860 45980
rect 206640 45860 206860 45910
rect 207140 46090 207360 46140
rect 207140 46020 207150 46090
rect 207350 46020 207360 46090
rect 207140 45980 207360 46020
rect 207140 45910 207150 45980
rect 207350 45910 207360 45980
rect 207140 45860 207360 45910
rect 207640 46090 207860 46140
rect 207640 46020 207650 46090
rect 207850 46020 207860 46090
rect 207640 45980 207860 46020
rect 207640 45910 207650 45980
rect 207850 45910 207860 45980
rect 207640 45860 207860 45910
rect 204000 45850 208000 45860
rect 204000 45650 204020 45850
rect 204090 45650 204410 45850
rect 204480 45650 204520 45850
rect 204590 45650 204910 45850
rect 204980 45650 205020 45850
rect 205090 45650 205410 45850
rect 205480 45650 205520 45850
rect 205590 45650 205910 45850
rect 205980 45650 206020 45850
rect 206090 45650 206410 45850
rect 206480 45650 206520 45850
rect 206590 45650 206910 45850
rect 206980 45650 207020 45850
rect 207090 45650 207410 45850
rect 207480 45650 207520 45850
rect 207590 45650 207910 45850
rect 207980 45650 208000 45850
rect 204000 45640 208000 45650
rect 204140 45590 204360 45640
rect 204140 45520 204150 45590
rect 204350 45520 204360 45590
rect 204140 45480 204360 45520
rect 204140 45410 204150 45480
rect 204350 45410 204360 45480
rect 204140 45360 204360 45410
rect 204640 45590 204860 45640
rect 204640 45520 204650 45590
rect 204850 45520 204860 45590
rect 204640 45480 204860 45520
rect 204640 45410 204650 45480
rect 204850 45410 204860 45480
rect 204640 45360 204860 45410
rect 205140 45590 205360 45640
rect 205140 45520 205150 45590
rect 205350 45520 205360 45590
rect 205140 45480 205360 45520
rect 205140 45410 205150 45480
rect 205350 45410 205360 45480
rect 205140 45360 205360 45410
rect 205640 45590 205860 45640
rect 205640 45520 205650 45590
rect 205850 45520 205860 45590
rect 205640 45480 205860 45520
rect 205640 45410 205650 45480
rect 205850 45410 205860 45480
rect 205640 45360 205860 45410
rect 206140 45590 206360 45640
rect 206140 45520 206150 45590
rect 206350 45520 206360 45590
rect 206140 45480 206360 45520
rect 206140 45410 206150 45480
rect 206350 45410 206360 45480
rect 206140 45360 206360 45410
rect 206640 45590 206860 45640
rect 206640 45520 206650 45590
rect 206850 45520 206860 45590
rect 206640 45480 206860 45520
rect 206640 45410 206650 45480
rect 206850 45410 206860 45480
rect 206640 45360 206860 45410
rect 207140 45590 207360 45640
rect 207140 45520 207150 45590
rect 207350 45520 207360 45590
rect 207140 45480 207360 45520
rect 207140 45410 207150 45480
rect 207350 45410 207360 45480
rect 207140 45360 207360 45410
rect 207640 45590 207860 45640
rect 207640 45520 207650 45590
rect 207850 45520 207860 45590
rect 207640 45480 207860 45520
rect 207640 45410 207650 45480
rect 207850 45410 207860 45480
rect 207640 45360 207860 45410
rect 204000 45350 208000 45360
rect 204000 45150 204020 45350
rect 204090 45150 204410 45350
rect 204480 45150 204520 45350
rect 204590 45150 204910 45350
rect 204980 45150 205020 45350
rect 205090 45150 205410 45350
rect 205480 45150 205520 45350
rect 205590 45150 205910 45350
rect 205980 45150 206020 45350
rect 206090 45150 206410 45350
rect 206480 45150 206520 45350
rect 206590 45150 206910 45350
rect 206980 45150 207020 45350
rect 207090 45150 207410 45350
rect 207480 45150 207520 45350
rect 207590 45150 207910 45350
rect 207980 45150 208000 45350
rect 204000 45140 208000 45150
rect 204140 45090 204360 45140
rect 204140 45020 204150 45090
rect 204350 45020 204360 45090
rect 204140 44980 204360 45020
rect 204140 44910 204150 44980
rect 204350 44910 204360 44980
rect 204140 44860 204360 44910
rect 204640 45090 204860 45140
rect 204640 45020 204650 45090
rect 204850 45020 204860 45090
rect 204640 44980 204860 45020
rect 204640 44910 204650 44980
rect 204850 44910 204860 44980
rect 204640 44860 204860 44910
rect 205140 45090 205360 45140
rect 205140 45020 205150 45090
rect 205350 45020 205360 45090
rect 205140 44980 205360 45020
rect 205140 44910 205150 44980
rect 205350 44910 205360 44980
rect 205140 44860 205360 44910
rect 205640 45090 205860 45140
rect 205640 45020 205650 45090
rect 205850 45020 205860 45090
rect 205640 44980 205860 45020
rect 205640 44910 205650 44980
rect 205850 44910 205860 44980
rect 205640 44860 205860 44910
rect 206140 45090 206360 45140
rect 206140 45020 206150 45090
rect 206350 45020 206360 45090
rect 206140 44980 206360 45020
rect 206140 44910 206150 44980
rect 206350 44910 206360 44980
rect 206140 44860 206360 44910
rect 206640 45090 206860 45140
rect 206640 45020 206650 45090
rect 206850 45020 206860 45090
rect 206640 44980 206860 45020
rect 206640 44910 206650 44980
rect 206850 44910 206860 44980
rect 206640 44860 206860 44910
rect 207140 45090 207360 45140
rect 207140 45020 207150 45090
rect 207350 45020 207360 45090
rect 207140 44980 207360 45020
rect 207140 44910 207150 44980
rect 207350 44910 207360 44980
rect 207140 44860 207360 44910
rect 207640 45090 207860 45140
rect 207640 45020 207650 45090
rect 207850 45020 207860 45090
rect 207640 44980 207860 45020
rect 207640 44910 207650 44980
rect 207850 44910 207860 44980
rect 207640 44860 207860 44910
rect 204000 44850 208000 44860
rect 204000 44650 204020 44850
rect 204090 44650 204410 44850
rect 204480 44650 204520 44850
rect 204590 44650 204910 44850
rect 204980 44650 205020 44850
rect 205090 44650 205410 44850
rect 205480 44650 205520 44850
rect 205590 44650 205910 44850
rect 205980 44650 206020 44850
rect 206090 44650 206410 44850
rect 206480 44650 206520 44850
rect 206590 44650 206910 44850
rect 206980 44650 207020 44850
rect 207090 44650 207410 44850
rect 207480 44650 207520 44850
rect 207590 44650 207910 44850
rect 207980 44650 208000 44850
rect 204000 44640 208000 44650
rect 204140 44590 204360 44640
rect 204140 44520 204150 44590
rect 204350 44520 204360 44590
rect 204140 44480 204360 44520
rect 204140 44410 204150 44480
rect 204350 44410 204360 44480
rect 204140 44360 204360 44410
rect 204640 44590 204860 44640
rect 204640 44520 204650 44590
rect 204850 44520 204860 44590
rect 204640 44480 204860 44520
rect 204640 44410 204650 44480
rect 204850 44410 204860 44480
rect 204640 44360 204860 44410
rect 205140 44590 205360 44640
rect 205140 44520 205150 44590
rect 205350 44520 205360 44590
rect 205140 44480 205360 44520
rect 205140 44410 205150 44480
rect 205350 44410 205360 44480
rect 205140 44360 205360 44410
rect 205640 44590 205860 44640
rect 205640 44520 205650 44590
rect 205850 44520 205860 44590
rect 205640 44480 205860 44520
rect 205640 44410 205650 44480
rect 205850 44410 205860 44480
rect 205640 44360 205860 44410
rect 206140 44590 206360 44640
rect 206140 44520 206150 44590
rect 206350 44520 206360 44590
rect 206140 44480 206360 44520
rect 206140 44410 206150 44480
rect 206350 44410 206360 44480
rect 206140 44360 206360 44410
rect 206640 44590 206860 44640
rect 206640 44520 206650 44590
rect 206850 44520 206860 44590
rect 206640 44480 206860 44520
rect 206640 44410 206650 44480
rect 206850 44410 206860 44480
rect 206640 44360 206860 44410
rect 207140 44590 207360 44640
rect 207140 44520 207150 44590
rect 207350 44520 207360 44590
rect 207140 44480 207360 44520
rect 207140 44410 207150 44480
rect 207350 44410 207360 44480
rect 207140 44360 207360 44410
rect 207640 44590 207860 44640
rect 207640 44520 207650 44590
rect 207850 44520 207860 44590
rect 207640 44480 207860 44520
rect 207640 44410 207650 44480
rect 207850 44410 207860 44480
rect 207640 44360 207860 44410
rect 204000 44350 208000 44360
rect 204000 44150 204020 44350
rect 204090 44150 204410 44350
rect 204480 44150 204520 44350
rect 204590 44150 204910 44350
rect 204980 44150 205020 44350
rect 205090 44150 205410 44350
rect 205480 44150 205520 44350
rect 205590 44150 205910 44350
rect 205980 44150 206020 44350
rect 206090 44150 206410 44350
rect 206480 44150 206520 44350
rect 206590 44150 206910 44350
rect 206980 44150 207020 44350
rect 207090 44150 207410 44350
rect 207480 44150 207520 44350
rect 207590 44150 207910 44350
rect 207980 44150 208000 44350
rect 204000 44140 208000 44150
rect 204140 44090 204360 44140
rect 204140 44020 204150 44090
rect 204350 44020 204360 44090
rect 204140 43980 204360 44020
rect 204140 43910 204150 43980
rect 204350 43910 204360 43980
rect 204140 43860 204360 43910
rect 204640 44090 204860 44140
rect 204640 44020 204650 44090
rect 204850 44020 204860 44090
rect 204640 43980 204860 44020
rect 204640 43910 204650 43980
rect 204850 43910 204860 43980
rect 204640 43860 204860 43910
rect 205140 44090 205360 44140
rect 205140 44020 205150 44090
rect 205350 44020 205360 44090
rect 205140 43980 205360 44020
rect 205140 43910 205150 43980
rect 205350 43910 205360 43980
rect 205140 43860 205360 43910
rect 205640 44090 205860 44140
rect 205640 44020 205650 44090
rect 205850 44020 205860 44090
rect 205640 43980 205860 44020
rect 205640 43910 205650 43980
rect 205850 43910 205860 43980
rect 205640 43860 205860 43910
rect 206140 44090 206360 44140
rect 206140 44020 206150 44090
rect 206350 44020 206360 44090
rect 206140 43980 206360 44020
rect 206140 43910 206150 43980
rect 206350 43910 206360 43980
rect 206140 43860 206360 43910
rect 206640 44090 206860 44140
rect 206640 44020 206650 44090
rect 206850 44020 206860 44090
rect 206640 43980 206860 44020
rect 206640 43910 206650 43980
rect 206850 43910 206860 43980
rect 206640 43860 206860 43910
rect 207140 44090 207360 44140
rect 207140 44020 207150 44090
rect 207350 44020 207360 44090
rect 207140 43980 207360 44020
rect 207140 43910 207150 43980
rect 207350 43910 207360 43980
rect 207140 43860 207360 43910
rect 207640 44090 207860 44140
rect 207640 44020 207650 44090
rect 207850 44020 207860 44090
rect 207640 43980 207860 44020
rect 207640 43910 207650 43980
rect 207850 43910 207860 43980
rect 207640 43860 207860 43910
rect 204000 43850 208000 43860
rect 204000 43650 204020 43850
rect 204090 43650 204410 43850
rect 204480 43650 204520 43850
rect 204590 43650 204910 43850
rect 204980 43650 205020 43850
rect 205090 43650 205410 43850
rect 205480 43650 205520 43850
rect 205590 43650 205910 43850
rect 205980 43650 206020 43850
rect 206090 43650 206410 43850
rect 206480 43650 206520 43850
rect 206590 43650 206910 43850
rect 206980 43650 207020 43850
rect 207090 43650 207410 43850
rect 207480 43650 207520 43850
rect 207590 43650 207910 43850
rect 207980 43650 208000 43850
rect 204000 43640 208000 43650
rect 204140 43590 204360 43640
rect 204140 43520 204150 43590
rect 204350 43520 204360 43590
rect 204140 43480 204360 43520
rect 204140 43410 204150 43480
rect 204350 43410 204360 43480
rect 204140 43360 204360 43410
rect 204640 43590 204860 43640
rect 204640 43520 204650 43590
rect 204850 43520 204860 43590
rect 204640 43480 204860 43520
rect 204640 43410 204650 43480
rect 204850 43410 204860 43480
rect 204640 43360 204860 43410
rect 205140 43590 205360 43640
rect 205140 43520 205150 43590
rect 205350 43520 205360 43590
rect 205140 43480 205360 43520
rect 205140 43410 205150 43480
rect 205350 43410 205360 43480
rect 205140 43360 205360 43410
rect 205640 43590 205860 43640
rect 205640 43520 205650 43590
rect 205850 43520 205860 43590
rect 205640 43480 205860 43520
rect 205640 43410 205650 43480
rect 205850 43410 205860 43480
rect 205640 43360 205860 43410
rect 206140 43590 206360 43640
rect 206140 43520 206150 43590
rect 206350 43520 206360 43590
rect 206140 43480 206360 43520
rect 206140 43410 206150 43480
rect 206350 43410 206360 43480
rect 206140 43360 206360 43410
rect 206640 43590 206860 43640
rect 206640 43520 206650 43590
rect 206850 43520 206860 43590
rect 206640 43480 206860 43520
rect 206640 43410 206650 43480
rect 206850 43410 206860 43480
rect 206640 43360 206860 43410
rect 207140 43590 207360 43640
rect 207140 43520 207150 43590
rect 207350 43520 207360 43590
rect 207140 43480 207360 43520
rect 207140 43410 207150 43480
rect 207350 43410 207360 43480
rect 207140 43360 207360 43410
rect 207640 43590 207860 43640
rect 207640 43520 207650 43590
rect 207850 43520 207860 43590
rect 207640 43480 207860 43520
rect 207640 43410 207650 43480
rect 207850 43410 207860 43480
rect 207640 43360 207860 43410
rect 204000 43350 208000 43360
rect 204000 43150 204020 43350
rect 204090 43150 204410 43350
rect 204480 43150 204520 43350
rect 204590 43150 204910 43350
rect 204980 43150 205020 43350
rect 205090 43150 205410 43350
rect 205480 43150 205520 43350
rect 205590 43150 205910 43350
rect 205980 43150 206020 43350
rect 206090 43150 206410 43350
rect 206480 43150 206520 43350
rect 206590 43150 206910 43350
rect 206980 43150 207020 43350
rect 207090 43150 207410 43350
rect 207480 43150 207520 43350
rect 207590 43150 207910 43350
rect 207980 43150 208000 43350
rect 204000 43140 208000 43150
rect 204140 43090 204360 43140
rect 204140 43020 204150 43090
rect 204350 43020 204360 43090
rect 204140 42980 204360 43020
rect 204140 42910 204150 42980
rect 204350 42910 204360 42980
rect 204140 42860 204360 42910
rect 204640 43090 204860 43140
rect 204640 43020 204650 43090
rect 204850 43020 204860 43090
rect 204640 42980 204860 43020
rect 204640 42910 204650 42980
rect 204850 42910 204860 42980
rect 204640 42860 204860 42910
rect 205140 43090 205360 43140
rect 205140 43020 205150 43090
rect 205350 43020 205360 43090
rect 205140 42980 205360 43020
rect 205140 42910 205150 42980
rect 205350 42910 205360 42980
rect 205140 42860 205360 42910
rect 205640 43090 205860 43140
rect 205640 43020 205650 43090
rect 205850 43020 205860 43090
rect 205640 42980 205860 43020
rect 205640 42910 205650 42980
rect 205850 42910 205860 42980
rect 205640 42860 205860 42910
rect 206140 43090 206360 43140
rect 206140 43020 206150 43090
rect 206350 43020 206360 43090
rect 206140 42980 206360 43020
rect 206140 42910 206150 42980
rect 206350 42910 206360 42980
rect 206140 42860 206360 42910
rect 206640 43090 206860 43140
rect 206640 43020 206650 43090
rect 206850 43020 206860 43090
rect 206640 42980 206860 43020
rect 206640 42910 206650 42980
rect 206850 42910 206860 42980
rect 206640 42860 206860 42910
rect 207140 43090 207360 43140
rect 207140 43020 207150 43090
rect 207350 43020 207360 43090
rect 207140 42980 207360 43020
rect 207140 42910 207150 42980
rect 207350 42910 207360 42980
rect 207140 42860 207360 42910
rect 207640 43090 207860 43140
rect 207640 43020 207650 43090
rect 207850 43020 207860 43090
rect 207640 42980 207860 43020
rect 207640 42910 207650 42980
rect 207850 42910 207860 42980
rect 207640 42860 207860 42910
rect 204000 42850 208000 42860
rect 204000 42650 204020 42850
rect 204090 42650 204410 42850
rect 204480 42650 204520 42850
rect 204590 42650 204910 42850
rect 204980 42650 205020 42850
rect 205090 42650 205410 42850
rect 205480 42650 205520 42850
rect 205590 42650 205910 42850
rect 205980 42650 206020 42850
rect 206090 42650 206410 42850
rect 206480 42650 206520 42850
rect 206590 42650 206910 42850
rect 206980 42650 207020 42850
rect 207090 42650 207410 42850
rect 207480 42650 207520 42850
rect 207590 42650 207910 42850
rect 207980 42650 208000 42850
rect 204000 42640 208000 42650
rect 204140 42590 204360 42640
rect 204140 42520 204150 42590
rect 204350 42520 204360 42590
rect 204140 42480 204360 42520
rect 204140 42410 204150 42480
rect 204350 42410 204360 42480
rect 204140 42360 204360 42410
rect 204640 42590 204860 42640
rect 204640 42520 204650 42590
rect 204850 42520 204860 42590
rect 204640 42480 204860 42520
rect 204640 42410 204650 42480
rect 204850 42410 204860 42480
rect 204640 42360 204860 42410
rect 205140 42590 205360 42640
rect 205140 42520 205150 42590
rect 205350 42520 205360 42590
rect 205140 42480 205360 42520
rect 205140 42410 205150 42480
rect 205350 42410 205360 42480
rect 205140 42360 205360 42410
rect 205640 42590 205860 42640
rect 205640 42520 205650 42590
rect 205850 42520 205860 42590
rect 205640 42480 205860 42520
rect 205640 42410 205650 42480
rect 205850 42410 205860 42480
rect 205640 42360 205860 42410
rect 206140 42590 206360 42640
rect 206140 42520 206150 42590
rect 206350 42520 206360 42590
rect 206140 42480 206360 42520
rect 206140 42410 206150 42480
rect 206350 42410 206360 42480
rect 206140 42360 206360 42410
rect 206640 42590 206860 42640
rect 206640 42520 206650 42590
rect 206850 42520 206860 42590
rect 206640 42480 206860 42520
rect 206640 42410 206650 42480
rect 206850 42410 206860 42480
rect 206640 42360 206860 42410
rect 207140 42590 207360 42640
rect 207140 42520 207150 42590
rect 207350 42520 207360 42590
rect 207140 42480 207360 42520
rect 207140 42410 207150 42480
rect 207350 42410 207360 42480
rect 207140 42360 207360 42410
rect 207640 42590 207860 42640
rect 207640 42520 207650 42590
rect 207850 42520 207860 42590
rect 207640 42480 207860 42520
rect 207640 42410 207650 42480
rect 207850 42410 207860 42480
rect 207640 42360 207860 42410
rect 204000 42350 208000 42360
rect 204000 42150 204020 42350
rect 204090 42150 204410 42350
rect 204480 42150 204520 42350
rect 204590 42150 204910 42350
rect 204980 42150 205020 42350
rect 205090 42150 205410 42350
rect 205480 42150 205520 42350
rect 205590 42150 205910 42350
rect 205980 42150 206020 42350
rect 206090 42150 206410 42350
rect 206480 42150 206520 42350
rect 206590 42150 206910 42350
rect 206980 42150 207020 42350
rect 207090 42150 207410 42350
rect 207480 42150 207520 42350
rect 207590 42150 207910 42350
rect 207980 42150 208000 42350
rect 204000 42140 208000 42150
rect 204140 42090 204360 42140
rect 204140 42020 204150 42090
rect 204350 42020 204360 42090
rect 204140 41980 204360 42020
rect 204140 41910 204150 41980
rect 204350 41910 204360 41980
rect 204140 41860 204360 41910
rect 204640 42090 204860 42140
rect 204640 42020 204650 42090
rect 204850 42020 204860 42090
rect 204640 41980 204860 42020
rect 204640 41910 204650 41980
rect 204850 41910 204860 41980
rect 204640 41860 204860 41910
rect 205140 42090 205360 42140
rect 205140 42020 205150 42090
rect 205350 42020 205360 42090
rect 205140 41980 205360 42020
rect 205140 41910 205150 41980
rect 205350 41910 205360 41980
rect 205140 41860 205360 41910
rect 205640 42090 205860 42140
rect 205640 42020 205650 42090
rect 205850 42020 205860 42090
rect 205640 41980 205860 42020
rect 205640 41910 205650 41980
rect 205850 41910 205860 41980
rect 205640 41860 205860 41910
rect 206140 42090 206360 42140
rect 206140 42020 206150 42090
rect 206350 42020 206360 42090
rect 206140 41980 206360 42020
rect 206140 41910 206150 41980
rect 206350 41910 206360 41980
rect 206140 41860 206360 41910
rect 206640 42090 206860 42140
rect 206640 42020 206650 42090
rect 206850 42020 206860 42090
rect 206640 41980 206860 42020
rect 206640 41910 206650 41980
rect 206850 41910 206860 41980
rect 206640 41860 206860 41910
rect 207140 42090 207360 42140
rect 207140 42020 207150 42090
rect 207350 42020 207360 42090
rect 207140 41980 207360 42020
rect 207140 41910 207150 41980
rect 207350 41910 207360 41980
rect 207140 41860 207360 41910
rect 207640 42090 207860 42140
rect 207640 42020 207650 42090
rect 207850 42020 207860 42090
rect 207640 41980 207860 42020
rect 207640 41910 207650 41980
rect 207850 41910 207860 41980
rect 207640 41860 207860 41910
rect 204000 41850 208000 41860
rect 204000 41650 204020 41850
rect 204090 41650 204410 41850
rect 204480 41650 204520 41850
rect 204590 41650 204910 41850
rect 204980 41650 205020 41850
rect 205090 41650 205410 41850
rect 205480 41650 205520 41850
rect 205590 41650 205910 41850
rect 205980 41650 206020 41850
rect 206090 41650 206410 41850
rect 206480 41650 206520 41850
rect 206590 41650 206910 41850
rect 206980 41650 207020 41850
rect 207090 41650 207410 41850
rect 207480 41650 207520 41850
rect 207590 41650 207910 41850
rect 207980 41650 208000 41850
rect 204000 41640 208000 41650
rect 204140 41590 204360 41640
rect 204140 41520 204150 41590
rect 204350 41520 204360 41590
rect 204140 41480 204360 41520
rect 204140 41410 204150 41480
rect 204350 41410 204360 41480
rect 204140 41360 204360 41410
rect 204640 41590 204860 41640
rect 204640 41520 204650 41590
rect 204850 41520 204860 41590
rect 204640 41480 204860 41520
rect 204640 41410 204650 41480
rect 204850 41410 204860 41480
rect 204640 41360 204860 41410
rect 205140 41590 205360 41640
rect 205140 41520 205150 41590
rect 205350 41520 205360 41590
rect 205140 41480 205360 41520
rect 205140 41410 205150 41480
rect 205350 41410 205360 41480
rect 205140 41360 205360 41410
rect 205640 41590 205860 41640
rect 205640 41520 205650 41590
rect 205850 41520 205860 41590
rect 205640 41480 205860 41520
rect 205640 41410 205650 41480
rect 205850 41410 205860 41480
rect 205640 41360 205860 41410
rect 206140 41590 206360 41640
rect 206140 41520 206150 41590
rect 206350 41520 206360 41590
rect 206140 41480 206360 41520
rect 206140 41410 206150 41480
rect 206350 41410 206360 41480
rect 206140 41360 206360 41410
rect 206640 41590 206860 41640
rect 206640 41520 206650 41590
rect 206850 41520 206860 41590
rect 206640 41480 206860 41520
rect 206640 41410 206650 41480
rect 206850 41410 206860 41480
rect 206640 41360 206860 41410
rect 207140 41590 207360 41640
rect 207140 41520 207150 41590
rect 207350 41520 207360 41590
rect 207140 41480 207360 41520
rect 207140 41410 207150 41480
rect 207350 41410 207360 41480
rect 207140 41360 207360 41410
rect 207640 41590 207860 41640
rect 207640 41520 207650 41590
rect 207850 41520 207860 41590
rect 207640 41480 207860 41520
rect 207640 41410 207650 41480
rect 207850 41410 207860 41480
rect 207640 41360 207860 41410
rect 204000 41350 208000 41360
rect 204000 41150 204020 41350
rect 204090 41150 204410 41350
rect 204480 41150 204520 41350
rect 204590 41150 204910 41350
rect 204980 41150 205020 41350
rect 205090 41150 205410 41350
rect 205480 41150 205520 41350
rect 205590 41150 205910 41350
rect 205980 41150 206020 41350
rect 206090 41150 206410 41350
rect 206480 41150 206520 41350
rect 206590 41150 206910 41350
rect 206980 41150 207020 41350
rect 207090 41150 207410 41350
rect 207480 41150 207520 41350
rect 207590 41150 207910 41350
rect 207980 41150 208000 41350
rect 204000 41140 208000 41150
rect 204140 41090 204360 41140
rect 204140 41020 204150 41090
rect 204350 41020 204360 41090
rect 204140 40980 204360 41020
rect 204140 40910 204150 40980
rect 204350 40910 204360 40980
rect 204140 40860 204360 40910
rect 204640 41090 204860 41140
rect 204640 41020 204650 41090
rect 204850 41020 204860 41090
rect 204640 40980 204860 41020
rect 204640 40910 204650 40980
rect 204850 40910 204860 40980
rect 204640 40860 204860 40910
rect 205140 41090 205360 41140
rect 205140 41020 205150 41090
rect 205350 41020 205360 41090
rect 205140 40980 205360 41020
rect 205140 40910 205150 40980
rect 205350 40910 205360 40980
rect 205140 40860 205360 40910
rect 205640 41090 205860 41140
rect 205640 41020 205650 41090
rect 205850 41020 205860 41090
rect 205640 40980 205860 41020
rect 205640 40910 205650 40980
rect 205850 40910 205860 40980
rect 205640 40860 205860 40910
rect 206140 41090 206360 41140
rect 206140 41020 206150 41090
rect 206350 41020 206360 41090
rect 206140 40980 206360 41020
rect 206140 40910 206150 40980
rect 206350 40910 206360 40980
rect 206140 40860 206360 40910
rect 206640 41090 206860 41140
rect 206640 41020 206650 41090
rect 206850 41020 206860 41090
rect 206640 40980 206860 41020
rect 206640 40910 206650 40980
rect 206850 40910 206860 40980
rect 206640 40860 206860 40910
rect 207140 41090 207360 41140
rect 207140 41020 207150 41090
rect 207350 41020 207360 41090
rect 207140 40980 207360 41020
rect 207140 40910 207150 40980
rect 207350 40910 207360 40980
rect 207140 40860 207360 40910
rect 207640 41090 207860 41140
rect 207640 41020 207650 41090
rect 207850 41020 207860 41090
rect 207640 40980 207860 41020
rect 207640 40910 207650 40980
rect 207850 40910 207860 40980
rect 207640 40860 207860 40910
rect 204000 40850 208000 40860
rect 204000 40650 204020 40850
rect 204090 40650 204410 40850
rect 204480 40650 204520 40850
rect 204590 40650 204910 40850
rect 204980 40650 205020 40850
rect 205090 40650 205410 40850
rect 205480 40650 205520 40850
rect 205590 40650 205910 40850
rect 205980 40650 206020 40850
rect 206090 40650 206410 40850
rect 206480 40650 206520 40850
rect 206590 40650 206910 40850
rect 206980 40650 207020 40850
rect 207090 40650 207410 40850
rect 207480 40650 207520 40850
rect 207590 40650 207910 40850
rect 207980 40650 208000 40850
rect 204000 40640 208000 40650
rect 204140 40590 204360 40640
rect 204140 40520 204150 40590
rect 204350 40520 204360 40590
rect 204140 40480 204360 40520
rect 204140 40410 204150 40480
rect 204350 40410 204360 40480
rect 204140 40360 204360 40410
rect 204640 40590 204860 40640
rect 204640 40520 204650 40590
rect 204850 40520 204860 40590
rect 204640 40480 204860 40520
rect 204640 40410 204650 40480
rect 204850 40410 204860 40480
rect 204640 40360 204860 40410
rect 205140 40590 205360 40640
rect 205140 40520 205150 40590
rect 205350 40520 205360 40590
rect 205140 40480 205360 40520
rect 205140 40410 205150 40480
rect 205350 40410 205360 40480
rect 205140 40360 205360 40410
rect 205640 40590 205860 40640
rect 205640 40520 205650 40590
rect 205850 40520 205860 40590
rect 205640 40480 205860 40520
rect 205640 40410 205650 40480
rect 205850 40410 205860 40480
rect 205640 40360 205860 40410
rect 206140 40590 206360 40640
rect 206140 40520 206150 40590
rect 206350 40520 206360 40590
rect 206140 40480 206360 40520
rect 206140 40410 206150 40480
rect 206350 40410 206360 40480
rect 206140 40360 206360 40410
rect 206640 40590 206860 40640
rect 206640 40520 206650 40590
rect 206850 40520 206860 40590
rect 206640 40480 206860 40520
rect 206640 40410 206650 40480
rect 206850 40410 206860 40480
rect 206640 40360 206860 40410
rect 207140 40590 207360 40640
rect 207140 40520 207150 40590
rect 207350 40520 207360 40590
rect 207140 40480 207360 40520
rect 207140 40410 207150 40480
rect 207350 40410 207360 40480
rect 207140 40360 207360 40410
rect 207640 40590 207860 40640
rect 207640 40520 207650 40590
rect 207850 40520 207860 40590
rect 207640 40480 207860 40520
rect 207640 40410 207650 40480
rect 207850 40410 207860 40480
rect 207640 40360 207860 40410
rect 204000 40350 208000 40360
rect 204000 40150 204020 40350
rect 204090 40150 204410 40350
rect 204480 40150 204520 40350
rect 204590 40150 204910 40350
rect 204980 40150 205020 40350
rect 205090 40150 205410 40350
rect 205480 40150 205520 40350
rect 205590 40150 205910 40350
rect 205980 40150 206020 40350
rect 206090 40150 206410 40350
rect 206480 40150 206520 40350
rect 206590 40150 206910 40350
rect 206980 40150 207020 40350
rect 207090 40150 207410 40350
rect 207480 40150 207520 40350
rect 207590 40150 207910 40350
rect 207980 40150 208000 40350
rect 204000 40140 208000 40150
rect 204140 40090 204360 40140
rect 204140 40020 204150 40090
rect 204350 40020 204360 40090
rect 204140 39980 204360 40020
rect 204140 39910 204150 39980
rect 204350 39910 204360 39980
rect 204140 39860 204360 39910
rect 204640 40090 204860 40140
rect 204640 40020 204650 40090
rect 204850 40020 204860 40090
rect 204640 39980 204860 40020
rect 204640 39910 204650 39980
rect 204850 39910 204860 39980
rect 204640 39860 204860 39910
rect 205140 40090 205360 40140
rect 205140 40020 205150 40090
rect 205350 40020 205360 40090
rect 205140 39980 205360 40020
rect 205140 39910 205150 39980
rect 205350 39910 205360 39980
rect 205140 39860 205360 39910
rect 205640 40090 205860 40140
rect 205640 40020 205650 40090
rect 205850 40020 205860 40090
rect 205640 39980 205860 40020
rect 205640 39910 205650 39980
rect 205850 39910 205860 39980
rect 205640 39860 205860 39910
rect 206140 40090 206360 40140
rect 206140 40020 206150 40090
rect 206350 40020 206360 40090
rect 206140 39980 206360 40020
rect 206140 39910 206150 39980
rect 206350 39910 206360 39980
rect 206140 39860 206360 39910
rect 206640 40090 206860 40140
rect 206640 40020 206650 40090
rect 206850 40020 206860 40090
rect 206640 39980 206860 40020
rect 206640 39910 206650 39980
rect 206850 39910 206860 39980
rect 206640 39860 206860 39910
rect 207140 40090 207360 40140
rect 207140 40020 207150 40090
rect 207350 40020 207360 40090
rect 207140 39980 207360 40020
rect 207140 39910 207150 39980
rect 207350 39910 207360 39980
rect 207140 39860 207360 39910
rect 207640 40090 207860 40140
rect 207640 40020 207650 40090
rect 207850 40020 207860 40090
rect 207640 39980 207860 40020
rect 207640 39910 207650 39980
rect 207850 39910 207860 39980
rect 207640 39860 207860 39910
rect 204000 39850 208000 39860
rect 204000 39650 204020 39850
rect 204090 39650 204410 39850
rect 204480 39650 204520 39850
rect 204590 39650 204910 39850
rect 204980 39650 205020 39850
rect 205090 39650 205410 39850
rect 205480 39650 205520 39850
rect 205590 39650 205910 39850
rect 205980 39650 206020 39850
rect 206090 39650 206410 39850
rect 206480 39650 206520 39850
rect 206590 39650 206910 39850
rect 206980 39650 207020 39850
rect 207090 39650 207410 39850
rect 207480 39650 207520 39850
rect 207590 39650 207910 39850
rect 207980 39650 208000 39850
rect 204000 39640 208000 39650
rect 204140 39590 204360 39640
rect 204140 39520 204150 39590
rect 204350 39520 204360 39590
rect 204140 39480 204360 39520
rect 204140 39410 204150 39480
rect 204350 39410 204360 39480
rect 204140 39360 204360 39410
rect 204640 39590 204860 39640
rect 204640 39520 204650 39590
rect 204850 39520 204860 39590
rect 204640 39480 204860 39520
rect 204640 39410 204650 39480
rect 204850 39410 204860 39480
rect 204640 39360 204860 39410
rect 205140 39590 205360 39640
rect 205140 39520 205150 39590
rect 205350 39520 205360 39590
rect 205140 39480 205360 39520
rect 205140 39410 205150 39480
rect 205350 39410 205360 39480
rect 205140 39360 205360 39410
rect 205640 39590 205860 39640
rect 205640 39520 205650 39590
rect 205850 39520 205860 39590
rect 205640 39480 205860 39520
rect 205640 39410 205650 39480
rect 205850 39410 205860 39480
rect 205640 39360 205860 39410
rect 206140 39590 206360 39640
rect 206140 39520 206150 39590
rect 206350 39520 206360 39590
rect 206140 39480 206360 39520
rect 206140 39410 206150 39480
rect 206350 39410 206360 39480
rect 206140 39360 206360 39410
rect 206640 39590 206860 39640
rect 206640 39520 206650 39590
rect 206850 39520 206860 39590
rect 206640 39480 206860 39520
rect 206640 39410 206650 39480
rect 206850 39410 206860 39480
rect 206640 39360 206860 39410
rect 207140 39590 207360 39640
rect 207140 39520 207150 39590
rect 207350 39520 207360 39590
rect 207140 39480 207360 39520
rect 207140 39410 207150 39480
rect 207350 39410 207360 39480
rect 207140 39360 207360 39410
rect 207640 39590 207860 39640
rect 207640 39520 207650 39590
rect 207850 39520 207860 39590
rect 207640 39480 207860 39520
rect 207640 39410 207650 39480
rect 207850 39410 207860 39480
rect 207640 39360 207860 39410
rect 204000 39350 208000 39360
rect 204000 39150 204020 39350
rect 204090 39150 204410 39350
rect 204480 39150 204520 39350
rect 204590 39150 204910 39350
rect 204980 39150 205020 39350
rect 205090 39150 205410 39350
rect 205480 39150 205520 39350
rect 205590 39150 205910 39350
rect 205980 39150 206020 39350
rect 206090 39150 206410 39350
rect 206480 39150 206520 39350
rect 206590 39150 206910 39350
rect 206980 39150 207020 39350
rect 207090 39150 207410 39350
rect 207480 39150 207520 39350
rect 207590 39150 207910 39350
rect 207980 39150 208000 39350
rect 204000 39140 208000 39150
rect 204140 39090 204360 39140
rect 204140 39020 204150 39090
rect 204350 39020 204360 39090
rect 204140 38980 204360 39020
rect 204140 38910 204150 38980
rect 204350 38910 204360 38980
rect 204140 38860 204360 38910
rect 204640 39090 204860 39140
rect 204640 39020 204650 39090
rect 204850 39020 204860 39090
rect 204640 38980 204860 39020
rect 204640 38910 204650 38980
rect 204850 38910 204860 38980
rect 204640 38860 204860 38910
rect 205140 39090 205360 39140
rect 205140 39020 205150 39090
rect 205350 39020 205360 39090
rect 205140 38980 205360 39020
rect 205140 38910 205150 38980
rect 205350 38910 205360 38980
rect 205140 38860 205360 38910
rect 205640 39090 205860 39140
rect 205640 39020 205650 39090
rect 205850 39020 205860 39090
rect 205640 38980 205860 39020
rect 205640 38910 205650 38980
rect 205850 38910 205860 38980
rect 205640 38860 205860 38910
rect 206140 39090 206360 39140
rect 206140 39020 206150 39090
rect 206350 39020 206360 39090
rect 206140 38980 206360 39020
rect 206140 38910 206150 38980
rect 206350 38910 206360 38980
rect 206140 38860 206360 38910
rect 206640 39090 206860 39140
rect 206640 39020 206650 39090
rect 206850 39020 206860 39090
rect 206640 38980 206860 39020
rect 206640 38910 206650 38980
rect 206850 38910 206860 38980
rect 206640 38860 206860 38910
rect 207140 39090 207360 39140
rect 207140 39020 207150 39090
rect 207350 39020 207360 39090
rect 207140 38980 207360 39020
rect 207140 38910 207150 38980
rect 207350 38910 207360 38980
rect 207140 38860 207360 38910
rect 207640 39090 207860 39140
rect 207640 39020 207650 39090
rect 207850 39020 207860 39090
rect 207640 38980 207860 39020
rect 207640 38910 207650 38980
rect 207850 38910 207860 38980
rect 207640 38860 207860 38910
rect 204000 38850 208000 38860
rect 204000 38650 204020 38850
rect 204090 38650 204410 38850
rect 204480 38650 204520 38850
rect 204590 38650 204910 38850
rect 204980 38650 205020 38850
rect 205090 38650 205410 38850
rect 205480 38650 205520 38850
rect 205590 38650 205910 38850
rect 205980 38650 206020 38850
rect 206090 38650 206410 38850
rect 206480 38650 206520 38850
rect 206590 38650 206910 38850
rect 206980 38650 207020 38850
rect 207090 38650 207410 38850
rect 207480 38650 207520 38850
rect 207590 38650 207910 38850
rect 207980 38650 208000 38850
rect 204000 38640 208000 38650
rect 204140 38590 204360 38640
rect 204140 38520 204150 38590
rect 204350 38520 204360 38590
rect 204140 38480 204360 38520
rect 204140 38410 204150 38480
rect 204350 38410 204360 38480
rect 204140 38360 204360 38410
rect 204640 38590 204860 38640
rect 204640 38520 204650 38590
rect 204850 38520 204860 38590
rect 204640 38480 204860 38520
rect 204640 38410 204650 38480
rect 204850 38410 204860 38480
rect 204640 38360 204860 38410
rect 205140 38590 205360 38640
rect 205140 38520 205150 38590
rect 205350 38520 205360 38590
rect 205140 38480 205360 38520
rect 205140 38410 205150 38480
rect 205350 38410 205360 38480
rect 205140 38360 205360 38410
rect 205640 38590 205860 38640
rect 205640 38520 205650 38590
rect 205850 38520 205860 38590
rect 205640 38480 205860 38520
rect 205640 38410 205650 38480
rect 205850 38410 205860 38480
rect 205640 38360 205860 38410
rect 206140 38590 206360 38640
rect 206140 38520 206150 38590
rect 206350 38520 206360 38590
rect 206140 38480 206360 38520
rect 206140 38410 206150 38480
rect 206350 38410 206360 38480
rect 206140 38360 206360 38410
rect 206640 38590 206860 38640
rect 206640 38520 206650 38590
rect 206850 38520 206860 38590
rect 206640 38480 206860 38520
rect 206640 38410 206650 38480
rect 206850 38410 206860 38480
rect 206640 38360 206860 38410
rect 207140 38590 207360 38640
rect 207140 38520 207150 38590
rect 207350 38520 207360 38590
rect 207140 38480 207360 38520
rect 207140 38410 207150 38480
rect 207350 38410 207360 38480
rect 207140 38360 207360 38410
rect 207640 38590 207860 38640
rect 207640 38520 207650 38590
rect 207850 38520 207860 38590
rect 207640 38480 207860 38520
rect 207640 38410 207650 38480
rect 207850 38410 207860 38480
rect 207640 38360 207860 38410
rect 204000 38350 208000 38360
rect 204000 38150 204020 38350
rect 204090 38150 204410 38350
rect 204480 38150 204520 38350
rect 204590 38150 204910 38350
rect 204980 38150 205020 38350
rect 205090 38150 205410 38350
rect 205480 38150 205520 38350
rect 205590 38150 205910 38350
rect 205980 38150 206020 38350
rect 206090 38150 206410 38350
rect 206480 38150 206520 38350
rect 206590 38150 206910 38350
rect 206980 38150 207020 38350
rect 207090 38150 207410 38350
rect 207480 38150 207520 38350
rect 207590 38150 207910 38350
rect 207980 38150 208000 38350
rect 204000 38140 208000 38150
rect 204140 38090 204360 38140
rect 204140 38020 204150 38090
rect 204350 38020 204360 38090
rect 204140 37980 204360 38020
rect 204140 37910 204150 37980
rect 204350 37910 204360 37980
rect 204140 37860 204360 37910
rect 204640 38090 204860 38140
rect 204640 38020 204650 38090
rect 204850 38020 204860 38090
rect 204640 37980 204860 38020
rect 204640 37910 204650 37980
rect 204850 37910 204860 37980
rect 204640 37860 204860 37910
rect 205140 38090 205360 38140
rect 205140 38020 205150 38090
rect 205350 38020 205360 38090
rect 205140 37980 205360 38020
rect 205140 37910 205150 37980
rect 205350 37910 205360 37980
rect 205140 37860 205360 37910
rect 205640 38090 205860 38140
rect 205640 38020 205650 38090
rect 205850 38020 205860 38090
rect 205640 37980 205860 38020
rect 205640 37910 205650 37980
rect 205850 37910 205860 37980
rect 205640 37860 205860 37910
rect 206140 38090 206360 38140
rect 206140 38020 206150 38090
rect 206350 38020 206360 38090
rect 206140 37980 206360 38020
rect 206140 37910 206150 37980
rect 206350 37910 206360 37980
rect 206140 37860 206360 37910
rect 206640 38090 206860 38140
rect 206640 38020 206650 38090
rect 206850 38020 206860 38090
rect 206640 37980 206860 38020
rect 206640 37910 206650 37980
rect 206850 37910 206860 37980
rect 206640 37860 206860 37910
rect 207140 38090 207360 38140
rect 207140 38020 207150 38090
rect 207350 38020 207360 38090
rect 207140 37980 207360 38020
rect 207140 37910 207150 37980
rect 207350 37910 207360 37980
rect 207140 37860 207360 37910
rect 207640 38090 207860 38140
rect 207640 38020 207650 38090
rect 207850 38020 207860 38090
rect 207640 37980 207860 38020
rect 207640 37910 207650 37980
rect 207850 37910 207860 37980
rect 207640 37860 207860 37910
rect 204000 37850 208000 37860
rect 204000 37650 204020 37850
rect 204090 37650 204410 37850
rect 204480 37650 204520 37850
rect 204590 37650 204910 37850
rect 204980 37650 205020 37850
rect 205090 37650 205410 37850
rect 205480 37650 205520 37850
rect 205590 37650 205910 37850
rect 205980 37650 206020 37850
rect 206090 37650 206410 37850
rect 206480 37650 206520 37850
rect 206590 37650 206910 37850
rect 206980 37650 207020 37850
rect 207090 37650 207410 37850
rect 207480 37650 207520 37850
rect 207590 37650 207910 37850
rect 207980 37650 208000 37850
rect 204000 37640 208000 37650
rect 204140 37590 204360 37640
rect 204140 37520 204150 37590
rect 204350 37520 204360 37590
rect 204140 37480 204360 37520
rect 204140 37410 204150 37480
rect 204350 37410 204360 37480
rect 204140 37360 204360 37410
rect 204640 37590 204860 37640
rect 204640 37520 204650 37590
rect 204850 37520 204860 37590
rect 204640 37480 204860 37520
rect 204640 37410 204650 37480
rect 204850 37410 204860 37480
rect 204640 37360 204860 37410
rect 205140 37590 205360 37640
rect 205140 37520 205150 37590
rect 205350 37520 205360 37590
rect 205140 37480 205360 37520
rect 205140 37410 205150 37480
rect 205350 37410 205360 37480
rect 205140 37360 205360 37410
rect 205640 37590 205860 37640
rect 205640 37520 205650 37590
rect 205850 37520 205860 37590
rect 205640 37480 205860 37520
rect 205640 37410 205650 37480
rect 205850 37410 205860 37480
rect 205640 37360 205860 37410
rect 206140 37590 206360 37640
rect 206140 37520 206150 37590
rect 206350 37520 206360 37590
rect 206140 37480 206360 37520
rect 206140 37410 206150 37480
rect 206350 37410 206360 37480
rect 206140 37360 206360 37410
rect 206640 37590 206860 37640
rect 206640 37520 206650 37590
rect 206850 37520 206860 37590
rect 206640 37480 206860 37520
rect 206640 37410 206650 37480
rect 206850 37410 206860 37480
rect 206640 37360 206860 37410
rect 207140 37590 207360 37640
rect 207140 37520 207150 37590
rect 207350 37520 207360 37590
rect 207140 37480 207360 37520
rect 207140 37410 207150 37480
rect 207350 37410 207360 37480
rect 207140 37360 207360 37410
rect 207640 37590 207860 37640
rect 207640 37520 207650 37590
rect 207850 37520 207860 37590
rect 207640 37480 207860 37520
rect 207640 37410 207650 37480
rect 207850 37410 207860 37480
rect 207640 37360 207860 37410
rect 204000 37350 208000 37360
rect 204000 37150 204020 37350
rect 204090 37150 204410 37350
rect 204480 37150 204520 37350
rect 204590 37150 204910 37350
rect 204980 37150 205020 37350
rect 205090 37150 205410 37350
rect 205480 37150 205520 37350
rect 205590 37150 205910 37350
rect 205980 37150 206020 37350
rect 206090 37150 206410 37350
rect 206480 37150 206520 37350
rect 206590 37150 206910 37350
rect 206980 37150 207020 37350
rect 207090 37150 207410 37350
rect 207480 37150 207520 37350
rect 207590 37150 207910 37350
rect 207980 37150 208000 37350
rect 204000 37140 208000 37150
rect 204140 37090 204360 37140
rect 204140 37020 204150 37090
rect 204350 37020 204360 37090
rect 204140 36980 204360 37020
rect 204140 36910 204150 36980
rect 204350 36910 204360 36980
rect 204140 36860 204360 36910
rect 204640 37090 204860 37140
rect 204640 37020 204650 37090
rect 204850 37020 204860 37090
rect 204640 36980 204860 37020
rect 204640 36910 204650 36980
rect 204850 36910 204860 36980
rect 204640 36860 204860 36910
rect 205140 37090 205360 37140
rect 205140 37020 205150 37090
rect 205350 37020 205360 37090
rect 205140 36980 205360 37020
rect 205140 36910 205150 36980
rect 205350 36910 205360 36980
rect 205140 36860 205360 36910
rect 205640 37090 205860 37140
rect 205640 37020 205650 37090
rect 205850 37020 205860 37090
rect 205640 36980 205860 37020
rect 205640 36910 205650 36980
rect 205850 36910 205860 36980
rect 205640 36860 205860 36910
rect 206140 37090 206360 37140
rect 206140 37020 206150 37090
rect 206350 37020 206360 37090
rect 206140 36980 206360 37020
rect 206140 36910 206150 36980
rect 206350 36910 206360 36980
rect 206140 36860 206360 36910
rect 206640 37090 206860 37140
rect 206640 37020 206650 37090
rect 206850 37020 206860 37090
rect 206640 36980 206860 37020
rect 206640 36910 206650 36980
rect 206850 36910 206860 36980
rect 206640 36860 206860 36910
rect 207140 37090 207360 37140
rect 207140 37020 207150 37090
rect 207350 37020 207360 37090
rect 207140 36980 207360 37020
rect 207140 36910 207150 36980
rect 207350 36910 207360 36980
rect 207140 36860 207360 36910
rect 207640 37090 207860 37140
rect 207640 37020 207650 37090
rect 207850 37020 207860 37090
rect 207640 36980 207860 37020
rect 207640 36910 207650 36980
rect 207850 36910 207860 36980
rect 207640 36860 207860 36910
rect 204000 36850 208000 36860
rect 204000 36650 204020 36850
rect 204090 36650 204410 36850
rect 204480 36650 204520 36850
rect 204590 36650 204910 36850
rect 204980 36650 205020 36850
rect 205090 36650 205410 36850
rect 205480 36650 205520 36850
rect 205590 36650 205910 36850
rect 205980 36650 206020 36850
rect 206090 36650 206410 36850
rect 206480 36650 206520 36850
rect 206590 36650 206910 36850
rect 206980 36650 207020 36850
rect 207090 36650 207410 36850
rect 207480 36650 207520 36850
rect 207590 36650 207910 36850
rect 207980 36650 208000 36850
rect 204000 36640 208000 36650
rect 204140 36590 204360 36640
rect 204140 36520 204150 36590
rect 204350 36520 204360 36590
rect 204140 36480 204360 36520
rect 204140 36410 204150 36480
rect 204350 36410 204360 36480
rect 204140 36360 204360 36410
rect 204640 36590 204860 36640
rect 204640 36520 204650 36590
rect 204850 36520 204860 36590
rect 204640 36480 204860 36520
rect 204640 36410 204650 36480
rect 204850 36410 204860 36480
rect 204640 36360 204860 36410
rect 205140 36590 205360 36640
rect 205140 36520 205150 36590
rect 205350 36520 205360 36590
rect 205140 36480 205360 36520
rect 205140 36410 205150 36480
rect 205350 36410 205360 36480
rect 205140 36360 205360 36410
rect 205640 36590 205860 36640
rect 205640 36520 205650 36590
rect 205850 36520 205860 36590
rect 205640 36480 205860 36520
rect 205640 36410 205650 36480
rect 205850 36410 205860 36480
rect 205640 36360 205860 36410
rect 206140 36590 206360 36640
rect 206140 36520 206150 36590
rect 206350 36520 206360 36590
rect 206140 36480 206360 36520
rect 206140 36410 206150 36480
rect 206350 36410 206360 36480
rect 206140 36360 206360 36410
rect 206640 36590 206860 36640
rect 206640 36520 206650 36590
rect 206850 36520 206860 36590
rect 206640 36480 206860 36520
rect 206640 36410 206650 36480
rect 206850 36410 206860 36480
rect 206640 36360 206860 36410
rect 207140 36590 207360 36640
rect 207140 36520 207150 36590
rect 207350 36520 207360 36590
rect 207140 36480 207360 36520
rect 207140 36410 207150 36480
rect 207350 36410 207360 36480
rect 207140 36360 207360 36410
rect 207640 36590 207860 36640
rect 207640 36520 207650 36590
rect 207850 36520 207860 36590
rect 207640 36480 207860 36520
rect 207640 36410 207650 36480
rect 207850 36410 207860 36480
rect 207640 36360 207860 36410
rect 204000 36350 208000 36360
rect 204000 36150 204020 36350
rect 204090 36150 204410 36350
rect 204480 36150 204520 36350
rect 204590 36150 204910 36350
rect 204980 36150 205020 36350
rect 205090 36150 205410 36350
rect 205480 36150 205520 36350
rect 205590 36150 205910 36350
rect 205980 36150 206020 36350
rect 206090 36150 206410 36350
rect 206480 36150 206520 36350
rect 206590 36150 206910 36350
rect 206980 36150 207020 36350
rect 207090 36150 207410 36350
rect 207480 36150 207520 36350
rect 207590 36150 207910 36350
rect 207980 36150 208000 36350
rect 204000 36140 208000 36150
rect 204140 36090 204360 36140
rect 204140 36020 204150 36090
rect 204350 36020 204360 36090
rect 204140 35980 204360 36020
rect 204140 35910 204150 35980
rect 204350 35910 204360 35980
rect 204140 35860 204360 35910
rect 204640 36090 204860 36140
rect 204640 36020 204650 36090
rect 204850 36020 204860 36090
rect 204640 35980 204860 36020
rect 204640 35910 204650 35980
rect 204850 35910 204860 35980
rect 204640 35860 204860 35910
rect 205140 36090 205360 36140
rect 205140 36020 205150 36090
rect 205350 36020 205360 36090
rect 205140 35980 205360 36020
rect 205140 35910 205150 35980
rect 205350 35910 205360 35980
rect 205140 35860 205360 35910
rect 205640 36090 205860 36140
rect 205640 36020 205650 36090
rect 205850 36020 205860 36090
rect 205640 35980 205860 36020
rect 205640 35910 205650 35980
rect 205850 35910 205860 35980
rect 205640 35860 205860 35910
rect 206140 36090 206360 36140
rect 206140 36020 206150 36090
rect 206350 36020 206360 36090
rect 206140 35980 206360 36020
rect 206140 35910 206150 35980
rect 206350 35910 206360 35980
rect 206140 35860 206360 35910
rect 206640 36090 206860 36140
rect 206640 36020 206650 36090
rect 206850 36020 206860 36090
rect 206640 35980 206860 36020
rect 206640 35910 206650 35980
rect 206850 35910 206860 35980
rect 206640 35860 206860 35910
rect 207140 36090 207360 36140
rect 207140 36020 207150 36090
rect 207350 36020 207360 36090
rect 207140 35980 207360 36020
rect 207140 35910 207150 35980
rect 207350 35910 207360 35980
rect 207140 35860 207360 35910
rect 207640 36090 207860 36140
rect 207640 36020 207650 36090
rect 207850 36020 207860 36090
rect 207640 35980 207860 36020
rect 207640 35910 207650 35980
rect 207850 35910 207860 35980
rect 207640 35860 207860 35910
rect 204000 35850 208000 35860
rect 204000 35650 204020 35850
rect 204090 35650 204410 35850
rect 204480 35650 204520 35850
rect 204590 35650 204910 35850
rect 204980 35650 205020 35850
rect 205090 35650 205410 35850
rect 205480 35650 205520 35850
rect 205590 35650 205910 35850
rect 205980 35650 206020 35850
rect 206090 35650 206410 35850
rect 206480 35650 206520 35850
rect 206590 35650 206910 35850
rect 206980 35650 207020 35850
rect 207090 35650 207410 35850
rect 207480 35650 207520 35850
rect 207590 35650 207910 35850
rect 207980 35650 208000 35850
rect 204000 35640 208000 35650
rect 204140 35590 204360 35640
rect 204140 35520 204150 35590
rect 204350 35520 204360 35590
rect 204140 35480 204360 35520
rect 204140 35410 204150 35480
rect 204350 35410 204360 35480
rect 204140 35360 204360 35410
rect 204640 35590 204860 35640
rect 204640 35520 204650 35590
rect 204850 35520 204860 35590
rect 204640 35480 204860 35520
rect 204640 35410 204650 35480
rect 204850 35410 204860 35480
rect 204640 35360 204860 35410
rect 205140 35590 205360 35640
rect 205140 35520 205150 35590
rect 205350 35520 205360 35590
rect 205140 35480 205360 35520
rect 205140 35410 205150 35480
rect 205350 35410 205360 35480
rect 205140 35360 205360 35410
rect 205640 35590 205860 35640
rect 205640 35520 205650 35590
rect 205850 35520 205860 35590
rect 205640 35480 205860 35520
rect 205640 35410 205650 35480
rect 205850 35410 205860 35480
rect 205640 35360 205860 35410
rect 206140 35590 206360 35640
rect 206140 35520 206150 35590
rect 206350 35520 206360 35590
rect 206140 35480 206360 35520
rect 206140 35410 206150 35480
rect 206350 35410 206360 35480
rect 206140 35360 206360 35410
rect 206640 35590 206860 35640
rect 206640 35520 206650 35590
rect 206850 35520 206860 35590
rect 206640 35480 206860 35520
rect 206640 35410 206650 35480
rect 206850 35410 206860 35480
rect 206640 35360 206860 35410
rect 207140 35590 207360 35640
rect 207140 35520 207150 35590
rect 207350 35520 207360 35590
rect 207140 35480 207360 35520
rect 207140 35410 207150 35480
rect 207350 35410 207360 35480
rect 207140 35360 207360 35410
rect 207640 35590 207860 35640
rect 207640 35520 207650 35590
rect 207850 35520 207860 35590
rect 207640 35480 207860 35520
rect 207640 35410 207650 35480
rect 207850 35410 207860 35480
rect 207640 35360 207860 35410
rect 204000 35350 208000 35360
rect 204000 35150 204020 35350
rect 204090 35150 204410 35350
rect 204480 35150 204520 35350
rect 204590 35150 204910 35350
rect 204980 35150 205020 35350
rect 205090 35150 205410 35350
rect 205480 35150 205520 35350
rect 205590 35150 205910 35350
rect 205980 35150 206020 35350
rect 206090 35150 206410 35350
rect 206480 35150 206520 35350
rect 206590 35150 206910 35350
rect 206980 35150 207020 35350
rect 207090 35150 207410 35350
rect 207480 35150 207520 35350
rect 207590 35150 207910 35350
rect 207980 35150 208000 35350
rect 204000 35140 208000 35150
rect 204140 35090 204360 35140
rect 204140 35020 204150 35090
rect 204350 35020 204360 35090
rect 204140 34980 204360 35020
rect 204140 34910 204150 34980
rect 204350 34910 204360 34980
rect 204140 34860 204360 34910
rect 204640 35090 204860 35140
rect 204640 35020 204650 35090
rect 204850 35020 204860 35090
rect 204640 34980 204860 35020
rect 204640 34910 204650 34980
rect 204850 34910 204860 34980
rect 204640 34860 204860 34910
rect 205140 35090 205360 35140
rect 205140 35020 205150 35090
rect 205350 35020 205360 35090
rect 205140 34980 205360 35020
rect 205140 34910 205150 34980
rect 205350 34910 205360 34980
rect 205140 34860 205360 34910
rect 205640 35090 205860 35140
rect 205640 35020 205650 35090
rect 205850 35020 205860 35090
rect 205640 34980 205860 35020
rect 205640 34910 205650 34980
rect 205850 34910 205860 34980
rect 205640 34860 205860 34910
rect 206140 35090 206360 35140
rect 206140 35020 206150 35090
rect 206350 35020 206360 35090
rect 206140 34980 206360 35020
rect 206140 34910 206150 34980
rect 206350 34910 206360 34980
rect 206140 34860 206360 34910
rect 206640 35090 206860 35140
rect 206640 35020 206650 35090
rect 206850 35020 206860 35090
rect 206640 34980 206860 35020
rect 206640 34910 206650 34980
rect 206850 34910 206860 34980
rect 206640 34860 206860 34910
rect 207140 35090 207360 35140
rect 207140 35020 207150 35090
rect 207350 35020 207360 35090
rect 207140 34980 207360 35020
rect 207140 34910 207150 34980
rect 207350 34910 207360 34980
rect 207140 34860 207360 34910
rect 207640 35090 207860 35140
rect 207640 35020 207650 35090
rect 207850 35020 207860 35090
rect 207640 34980 207860 35020
rect 207640 34910 207650 34980
rect 207850 34910 207860 34980
rect 207640 34860 207860 34910
rect 204000 34850 208000 34860
rect 204000 34650 204020 34850
rect 204090 34650 204410 34850
rect 204480 34650 204520 34850
rect 204590 34650 204910 34850
rect 204980 34650 205020 34850
rect 205090 34650 205410 34850
rect 205480 34650 205520 34850
rect 205590 34650 205910 34850
rect 205980 34650 206020 34850
rect 206090 34650 206410 34850
rect 206480 34650 206520 34850
rect 206590 34650 206910 34850
rect 206980 34650 207020 34850
rect 207090 34650 207410 34850
rect 207480 34650 207520 34850
rect 207590 34650 207910 34850
rect 207980 34650 208000 34850
rect 204000 34640 208000 34650
rect 204140 34590 204360 34640
rect 204140 34520 204150 34590
rect 204350 34520 204360 34590
rect 204140 34480 204360 34520
rect 204140 34410 204150 34480
rect 204350 34410 204360 34480
rect 204140 34360 204360 34410
rect 204640 34590 204860 34640
rect 204640 34520 204650 34590
rect 204850 34520 204860 34590
rect 204640 34480 204860 34520
rect 204640 34410 204650 34480
rect 204850 34410 204860 34480
rect 204640 34360 204860 34410
rect 205140 34590 205360 34640
rect 205140 34520 205150 34590
rect 205350 34520 205360 34590
rect 205140 34480 205360 34520
rect 205140 34410 205150 34480
rect 205350 34410 205360 34480
rect 205140 34360 205360 34410
rect 205640 34590 205860 34640
rect 205640 34520 205650 34590
rect 205850 34520 205860 34590
rect 205640 34480 205860 34520
rect 205640 34410 205650 34480
rect 205850 34410 205860 34480
rect 205640 34360 205860 34410
rect 206140 34590 206360 34640
rect 206140 34520 206150 34590
rect 206350 34520 206360 34590
rect 206140 34480 206360 34520
rect 206140 34410 206150 34480
rect 206350 34410 206360 34480
rect 206140 34360 206360 34410
rect 206640 34590 206860 34640
rect 206640 34520 206650 34590
rect 206850 34520 206860 34590
rect 206640 34480 206860 34520
rect 206640 34410 206650 34480
rect 206850 34410 206860 34480
rect 206640 34360 206860 34410
rect 207140 34590 207360 34640
rect 207140 34520 207150 34590
rect 207350 34520 207360 34590
rect 207140 34480 207360 34520
rect 207140 34410 207150 34480
rect 207350 34410 207360 34480
rect 207140 34360 207360 34410
rect 207640 34590 207860 34640
rect 207640 34520 207650 34590
rect 207850 34520 207860 34590
rect 207640 34480 207860 34520
rect 207640 34410 207650 34480
rect 207850 34410 207860 34480
rect 207640 34360 207860 34410
rect 204000 34350 208000 34360
rect 204000 34150 204020 34350
rect 204090 34150 204410 34350
rect 204480 34150 204520 34350
rect 204590 34150 204910 34350
rect 204980 34150 205020 34350
rect 205090 34150 205410 34350
rect 205480 34150 205520 34350
rect 205590 34150 205910 34350
rect 205980 34150 206020 34350
rect 206090 34150 206410 34350
rect 206480 34150 206520 34350
rect 206590 34150 206910 34350
rect 206980 34150 207020 34350
rect 207090 34150 207410 34350
rect 207480 34150 207520 34350
rect 207590 34150 207910 34350
rect 207980 34150 208000 34350
rect 204000 34140 208000 34150
rect 204140 34090 204360 34140
rect 204140 34020 204150 34090
rect 204350 34020 204360 34090
rect 204140 33980 204360 34020
rect 204140 33910 204150 33980
rect 204350 33910 204360 33980
rect 204140 33860 204360 33910
rect 204640 34090 204860 34140
rect 204640 34020 204650 34090
rect 204850 34020 204860 34090
rect 204640 33980 204860 34020
rect 204640 33910 204650 33980
rect 204850 33910 204860 33980
rect 204640 33860 204860 33910
rect 205140 34090 205360 34140
rect 205140 34020 205150 34090
rect 205350 34020 205360 34090
rect 205140 33980 205360 34020
rect 205140 33910 205150 33980
rect 205350 33910 205360 33980
rect 205140 33860 205360 33910
rect 205640 34090 205860 34140
rect 205640 34020 205650 34090
rect 205850 34020 205860 34090
rect 205640 33980 205860 34020
rect 205640 33910 205650 33980
rect 205850 33910 205860 33980
rect 205640 33860 205860 33910
rect 206140 34090 206360 34140
rect 206140 34020 206150 34090
rect 206350 34020 206360 34090
rect 206140 33980 206360 34020
rect 206140 33910 206150 33980
rect 206350 33910 206360 33980
rect 206140 33860 206360 33910
rect 206640 34090 206860 34140
rect 206640 34020 206650 34090
rect 206850 34020 206860 34090
rect 206640 33980 206860 34020
rect 206640 33910 206650 33980
rect 206850 33910 206860 33980
rect 206640 33860 206860 33910
rect 207140 34090 207360 34140
rect 207140 34020 207150 34090
rect 207350 34020 207360 34090
rect 207140 33980 207360 34020
rect 207140 33910 207150 33980
rect 207350 33910 207360 33980
rect 207140 33860 207360 33910
rect 207640 34090 207860 34140
rect 207640 34020 207650 34090
rect 207850 34020 207860 34090
rect 207640 33980 207860 34020
rect 207640 33910 207650 33980
rect 207850 33910 207860 33980
rect 207640 33860 207860 33910
rect 204000 33850 208000 33860
rect 204000 33650 204020 33850
rect 204090 33650 204410 33850
rect 204480 33650 204520 33850
rect 204590 33650 204910 33850
rect 204980 33650 205020 33850
rect 205090 33650 205410 33850
rect 205480 33650 205520 33850
rect 205590 33650 205910 33850
rect 205980 33650 206020 33850
rect 206090 33650 206410 33850
rect 206480 33650 206520 33850
rect 206590 33650 206910 33850
rect 206980 33650 207020 33850
rect 207090 33650 207410 33850
rect 207480 33650 207520 33850
rect 207590 33650 207910 33850
rect 207980 33650 208000 33850
rect 204000 33640 208000 33650
rect 204140 33590 204360 33640
rect 204140 33520 204150 33590
rect 204350 33520 204360 33590
rect 204140 33480 204360 33520
rect 204140 33410 204150 33480
rect 204350 33410 204360 33480
rect 204140 33360 204360 33410
rect 204640 33590 204860 33640
rect 204640 33520 204650 33590
rect 204850 33520 204860 33590
rect 204640 33480 204860 33520
rect 204640 33410 204650 33480
rect 204850 33410 204860 33480
rect 204640 33360 204860 33410
rect 205140 33590 205360 33640
rect 205140 33520 205150 33590
rect 205350 33520 205360 33590
rect 205140 33480 205360 33520
rect 205140 33410 205150 33480
rect 205350 33410 205360 33480
rect 205140 33360 205360 33410
rect 205640 33590 205860 33640
rect 205640 33520 205650 33590
rect 205850 33520 205860 33590
rect 205640 33480 205860 33520
rect 205640 33410 205650 33480
rect 205850 33410 205860 33480
rect 205640 33360 205860 33410
rect 206140 33590 206360 33640
rect 206140 33520 206150 33590
rect 206350 33520 206360 33590
rect 206140 33480 206360 33520
rect 206140 33410 206150 33480
rect 206350 33410 206360 33480
rect 206140 33360 206360 33410
rect 206640 33590 206860 33640
rect 206640 33520 206650 33590
rect 206850 33520 206860 33590
rect 206640 33480 206860 33520
rect 206640 33410 206650 33480
rect 206850 33410 206860 33480
rect 206640 33360 206860 33410
rect 207140 33590 207360 33640
rect 207140 33520 207150 33590
rect 207350 33520 207360 33590
rect 207140 33480 207360 33520
rect 207140 33410 207150 33480
rect 207350 33410 207360 33480
rect 207140 33360 207360 33410
rect 207640 33590 207860 33640
rect 207640 33520 207650 33590
rect 207850 33520 207860 33590
rect 207640 33480 207860 33520
rect 207640 33410 207650 33480
rect 207850 33410 207860 33480
rect 207640 33360 207860 33410
rect 204000 33350 208000 33360
rect 204000 33150 204020 33350
rect 204090 33150 204410 33350
rect 204480 33150 204520 33350
rect 204590 33150 204910 33350
rect 204980 33150 205020 33350
rect 205090 33150 205410 33350
rect 205480 33150 205520 33350
rect 205590 33150 205910 33350
rect 205980 33150 206020 33350
rect 206090 33150 206410 33350
rect 206480 33150 206520 33350
rect 206590 33150 206910 33350
rect 206980 33150 207020 33350
rect 207090 33150 207410 33350
rect 207480 33150 207520 33350
rect 207590 33150 207910 33350
rect 207980 33150 208000 33350
rect 204000 33140 208000 33150
rect 204140 33090 204360 33140
rect 204140 33020 204150 33090
rect 204350 33020 204360 33090
rect 204140 32980 204360 33020
rect 204140 32910 204150 32980
rect 204350 32910 204360 32980
rect 204140 32860 204360 32910
rect 204640 33090 204860 33140
rect 204640 33020 204650 33090
rect 204850 33020 204860 33090
rect 204640 32980 204860 33020
rect 204640 32910 204650 32980
rect 204850 32910 204860 32980
rect 204640 32860 204860 32910
rect 205140 33090 205360 33140
rect 205140 33020 205150 33090
rect 205350 33020 205360 33090
rect 205140 32980 205360 33020
rect 205140 32910 205150 32980
rect 205350 32910 205360 32980
rect 205140 32860 205360 32910
rect 205640 33090 205860 33140
rect 205640 33020 205650 33090
rect 205850 33020 205860 33090
rect 205640 32980 205860 33020
rect 205640 32910 205650 32980
rect 205850 32910 205860 32980
rect 205640 32860 205860 32910
rect 206140 33090 206360 33140
rect 206140 33020 206150 33090
rect 206350 33020 206360 33090
rect 206140 32980 206360 33020
rect 206140 32910 206150 32980
rect 206350 32910 206360 32980
rect 206140 32860 206360 32910
rect 206640 33090 206860 33140
rect 206640 33020 206650 33090
rect 206850 33020 206860 33090
rect 206640 32980 206860 33020
rect 206640 32910 206650 32980
rect 206850 32910 206860 32980
rect 206640 32860 206860 32910
rect 207140 33090 207360 33140
rect 207140 33020 207150 33090
rect 207350 33020 207360 33090
rect 207140 32980 207360 33020
rect 207140 32910 207150 32980
rect 207350 32910 207360 32980
rect 207140 32860 207360 32910
rect 207640 33090 207860 33140
rect 207640 33020 207650 33090
rect 207850 33020 207860 33090
rect 207640 32980 207860 33020
rect 207640 32910 207650 32980
rect 207850 32910 207860 32980
rect 207640 32860 207860 32910
rect 204000 32850 208000 32860
rect 204000 32650 204020 32850
rect 204090 32650 204410 32850
rect 204480 32650 204520 32850
rect 204590 32650 204910 32850
rect 204980 32650 205020 32850
rect 205090 32650 205410 32850
rect 205480 32650 205520 32850
rect 205590 32650 205910 32850
rect 205980 32650 206020 32850
rect 206090 32650 206410 32850
rect 206480 32650 206520 32850
rect 206590 32650 206910 32850
rect 206980 32650 207020 32850
rect 207090 32650 207410 32850
rect 207480 32650 207520 32850
rect 207590 32650 207910 32850
rect 207980 32650 208000 32850
rect 204000 32640 208000 32650
rect 204140 32590 204360 32640
rect 204140 32520 204150 32590
rect 204350 32520 204360 32590
rect 204140 32480 204360 32520
rect 204140 32410 204150 32480
rect 204350 32410 204360 32480
rect 204140 32360 204360 32410
rect 204640 32590 204860 32640
rect 204640 32520 204650 32590
rect 204850 32520 204860 32590
rect 204640 32480 204860 32520
rect 204640 32410 204650 32480
rect 204850 32410 204860 32480
rect 204640 32360 204860 32410
rect 205140 32590 205360 32640
rect 205140 32520 205150 32590
rect 205350 32520 205360 32590
rect 205140 32480 205360 32520
rect 205140 32410 205150 32480
rect 205350 32410 205360 32480
rect 205140 32360 205360 32410
rect 205640 32590 205860 32640
rect 205640 32520 205650 32590
rect 205850 32520 205860 32590
rect 205640 32480 205860 32520
rect 205640 32410 205650 32480
rect 205850 32410 205860 32480
rect 205640 32360 205860 32410
rect 206140 32590 206360 32640
rect 206140 32520 206150 32590
rect 206350 32520 206360 32590
rect 206140 32480 206360 32520
rect 206140 32410 206150 32480
rect 206350 32410 206360 32480
rect 206140 32360 206360 32410
rect 206640 32590 206860 32640
rect 206640 32520 206650 32590
rect 206850 32520 206860 32590
rect 206640 32480 206860 32520
rect 206640 32410 206650 32480
rect 206850 32410 206860 32480
rect 206640 32360 206860 32410
rect 207140 32590 207360 32640
rect 207140 32520 207150 32590
rect 207350 32520 207360 32590
rect 207140 32480 207360 32520
rect 207140 32410 207150 32480
rect 207350 32410 207360 32480
rect 207140 32360 207360 32410
rect 207640 32590 207860 32640
rect 207640 32520 207650 32590
rect 207850 32520 207860 32590
rect 207640 32480 207860 32520
rect 207640 32410 207650 32480
rect 207850 32410 207860 32480
rect 207640 32360 207860 32410
rect 204000 32350 208000 32360
rect 204000 32150 204020 32350
rect 204090 32150 204410 32350
rect 204480 32150 204520 32350
rect 204590 32150 204910 32350
rect 204980 32150 205020 32350
rect 205090 32150 205410 32350
rect 205480 32150 205520 32350
rect 205590 32150 205910 32350
rect 205980 32150 206020 32350
rect 206090 32150 206410 32350
rect 206480 32150 206520 32350
rect 206590 32150 206910 32350
rect 206980 32150 207020 32350
rect 207090 32150 207410 32350
rect 207480 32150 207520 32350
rect 207590 32150 207910 32350
rect 207980 32150 208000 32350
rect 204000 32140 208000 32150
rect 204140 32090 204360 32140
rect 204140 32020 204150 32090
rect 204350 32020 204360 32090
rect 204140 31980 204360 32020
rect 204140 31910 204150 31980
rect 204350 31910 204360 31980
rect 204140 31860 204360 31910
rect 204640 32090 204860 32140
rect 204640 32020 204650 32090
rect 204850 32020 204860 32090
rect 204640 31980 204860 32020
rect 204640 31910 204650 31980
rect 204850 31910 204860 31980
rect 204640 31860 204860 31910
rect 205140 32090 205360 32140
rect 205140 32020 205150 32090
rect 205350 32020 205360 32090
rect 205140 31980 205360 32020
rect 205140 31910 205150 31980
rect 205350 31910 205360 31980
rect 205140 31860 205360 31910
rect 205640 32090 205860 32140
rect 205640 32020 205650 32090
rect 205850 32020 205860 32090
rect 205640 31980 205860 32020
rect 205640 31910 205650 31980
rect 205850 31910 205860 31980
rect 205640 31860 205860 31910
rect 206140 32090 206360 32140
rect 206140 32020 206150 32090
rect 206350 32020 206360 32090
rect 206140 31980 206360 32020
rect 206140 31910 206150 31980
rect 206350 31910 206360 31980
rect 206140 31860 206360 31910
rect 206640 32090 206860 32140
rect 206640 32020 206650 32090
rect 206850 32020 206860 32090
rect 206640 31980 206860 32020
rect 206640 31910 206650 31980
rect 206850 31910 206860 31980
rect 206640 31860 206860 31910
rect 207140 32090 207360 32140
rect 207140 32020 207150 32090
rect 207350 32020 207360 32090
rect 207140 31980 207360 32020
rect 207140 31910 207150 31980
rect 207350 31910 207360 31980
rect 207140 31860 207360 31910
rect 207640 32090 207860 32140
rect 207640 32020 207650 32090
rect 207850 32020 207860 32090
rect 207640 31980 207860 32020
rect 207640 31910 207650 31980
rect 207850 31910 207860 31980
rect 207640 31860 207860 31910
rect 204000 31850 208000 31860
rect 204000 31650 204020 31850
rect 204090 31650 204410 31850
rect 204480 31650 204520 31850
rect 204590 31650 204910 31850
rect 204980 31650 205020 31850
rect 205090 31650 205410 31850
rect 205480 31650 205520 31850
rect 205590 31650 205910 31850
rect 205980 31650 206020 31850
rect 206090 31650 206410 31850
rect 206480 31650 206520 31850
rect 206590 31650 206910 31850
rect 206980 31650 207020 31850
rect 207090 31650 207410 31850
rect 207480 31650 207520 31850
rect 207590 31650 207910 31850
rect 207980 31650 208000 31850
rect 204000 31640 208000 31650
rect 204140 31590 204360 31640
rect 204140 31520 204150 31590
rect 204350 31520 204360 31590
rect 204140 31480 204360 31520
rect 204140 31410 204150 31480
rect 204350 31410 204360 31480
rect 204140 31360 204360 31410
rect 204640 31590 204860 31640
rect 204640 31520 204650 31590
rect 204850 31520 204860 31590
rect 204640 31480 204860 31520
rect 204640 31410 204650 31480
rect 204850 31410 204860 31480
rect 204640 31360 204860 31410
rect 205140 31590 205360 31640
rect 205140 31520 205150 31590
rect 205350 31520 205360 31590
rect 205140 31480 205360 31520
rect 205140 31410 205150 31480
rect 205350 31410 205360 31480
rect 205140 31360 205360 31410
rect 205640 31590 205860 31640
rect 205640 31520 205650 31590
rect 205850 31520 205860 31590
rect 205640 31480 205860 31520
rect 205640 31410 205650 31480
rect 205850 31410 205860 31480
rect 205640 31360 205860 31410
rect 206140 31590 206360 31640
rect 206140 31520 206150 31590
rect 206350 31520 206360 31590
rect 206140 31480 206360 31520
rect 206140 31410 206150 31480
rect 206350 31410 206360 31480
rect 206140 31360 206360 31410
rect 206640 31590 206860 31640
rect 206640 31520 206650 31590
rect 206850 31520 206860 31590
rect 206640 31480 206860 31520
rect 206640 31410 206650 31480
rect 206850 31410 206860 31480
rect 206640 31360 206860 31410
rect 207140 31590 207360 31640
rect 207140 31520 207150 31590
rect 207350 31520 207360 31590
rect 207140 31480 207360 31520
rect 207140 31410 207150 31480
rect 207350 31410 207360 31480
rect 207140 31360 207360 31410
rect 207640 31590 207860 31640
rect 207640 31520 207650 31590
rect 207850 31520 207860 31590
rect 207640 31480 207860 31520
rect 207640 31410 207650 31480
rect 207850 31410 207860 31480
rect 207640 31360 207860 31410
rect 204000 31350 208000 31360
rect 204000 31150 204020 31350
rect 204090 31150 204410 31350
rect 204480 31150 204520 31350
rect 204590 31150 204910 31350
rect 204980 31150 205020 31350
rect 205090 31150 205410 31350
rect 205480 31150 205520 31350
rect 205590 31150 205910 31350
rect 205980 31150 206020 31350
rect 206090 31150 206410 31350
rect 206480 31150 206520 31350
rect 206590 31150 206910 31350
rect 206980 31150 207020 31350
rect 207090 31150 207410 31350
rect 207480 31150 207520 31350
rect 207590 31150 207910 31350
rect 207980 31150 208000 31350
rect 204000 31140 208000 31150
rect 204140 31090 204360 31140
rect 204140 31020 204150 31090
rect 204350 31020 204360 31090
rect 204140 30980 204360 31020
rect 204140 30910 204150 30980
rect 204350 30910 204360 30980
rect 204140 30860 204360 30910
rect 204640 31090 204860 31140
rect 204640 31020 204650 31090
rect 204850 31020 204860 31090
rect 204640 30980 204860 31020
rect 204640 30910 204650 30980
rect 204850 30910 204860 30980
rect 204640 30860 204860 30910
rect 205140 31090 205360 31140
rect 205140 31020 205150 31090
rect 205350 31020 205360 31090
rect 205140 30980 205360 31020
rect 205140 30910 205150 30980
rect 205350 30910 205360 30980
rect 205140 30860 205360 30910
rect 205640 31090 205860 31140
rect 205640 31020 205650 31090
rect 205850 31020 205860 31090
rect 205640 30980 205860 31020
rect 205640 30910 205650 30980
rect 205850 30910 205860 30980
rect 205640 30860 205860 30910
rect 206140 31090 206360 31140
rect 206140 31020 206150 31090
rect 206350 31020 206360 31090
rect 206140 30980 206360 31020
rect 206140 30910 206150 30980
rect 206350 30910 206360 30980
rect 206140 30860 206360 30910
rect 206640 31090 206860 31140
rect 206640 31020 206650 31090
rect 206850 31020 206860 31090
rect 206640 30980 206860 31020
rect 206640 30910 206650 30980
rect 206850 30910 206860 30980
rect 206640 30860 206860 30910
rect 207140 31090 207360 31140
rect 207140 31020 207150 31090
rect 207350 31020 207360 31090
rect 207140 30980 207360 31020
rect 207140 30910 207150 30980
rect 207350 30910 207360 30980
rect 207140 30860 207360 30910
rect 207640 31090 207860 31140
rect 207640 31020 207650 31090
rect 207850 31020 207860 31090
rect 207640 30980 207860 31020
rect 207640 30910 207650 30980
rect 207850 30910 207860 30980
rect 207640 30860 207860 30910
rect 204000 30850 208000 30860
rect 204000 30650 204020 30850
rect 204090 30650 204410 30850
rect 204480 30650 204520 30850
rect 204590 30650 204910 30850
rect 204980 30650 205020 30850
rect 205090 30650 205410 30850
rect 205480 30650 205520 30850
rect 205590 30650 205910 30850
rect 205980 30650 206020 30850
rect 206090 30650 206410 30850
rect 206480 30650 206520 30850
rect 206590 30650 206910 30850
rect 206980 30650 207020 30850
rect 207090 30650 207410 30850
rect 207480 30650 207520 30850
rect 207590 30650 207910 30850
rect 207980 30650 208000 30850
rect 204000 30640 208000 30650
rect 204140 30590 204360 30640
rect 204140 30520 204150 30590
rect 204350 30520 204360 30590
rect 204140 30480 204360 30520
rect 204140 30410 204150 30480
rect 204350 30410 204360 30480
rect 204140 30360 204360 30410
rect 204640 30590 204860 30640
rect 204640 30520 204650 30590
rect 204850 30520 204860 30590
rect 204640 30480 204860 30520
rect 204640 30410 204650 30480
rect 204850 30410 204860 30480
rect 204640 30360 204860 30410
rect 205140 30590 205360 30640
rect 205140 30520 205150 30590
rect 205350 30520 205360 30590
rect 205140 30480 205360 30520
rect 205140 30410 205150 30480
rect 205350 30410 205360 30480
rect 205140 30360 205360 30410
rect 205640 30590 205860 30640
rect 205640 30520 205650 30590
rect 205850 30520 205860 30590
rect 205640 30480 205860 30520
rect 205640 30410 205650 30480
rect 205850 30410 205860 30480
rect 205640 30360 205860 30410
rect 206140 30590 206360 30640
rect 206140 30520 206150 30590
rect 206350 30520 206360 30590
rect 206140 30480 206360 30520
rect 206140 30410 206150 30480
rect 206350 30410 206360 30480
rect 206140 30360 206360 30410
rect 206640 30590 206860 30640
rect 206640 30520 206650 30590
rect 206850 30520 206860 30590
rect 206640 30480 206860 30520
rect 206640 30410 206650 30480
rect 206850 30410 206860 30480
rect 206640 30360 206860 30410
rect 207140 30590 207360 30640
rect 207140 30520 207150 30590
rect 207350 30520 207360 30590
rect 207140 30480 207360 30520
rect 207140 30410 207150 30480
rect 207350 30410 207360 30480
rect 207140 30360 207360 30410
rect 207640 30590 207860 30640
rect 207640 30520 207650 30590
rect 207850 30520 207860 30590
rect 207640 30480 207860 30520
rect 207640 30410 207650 30480
rect 207850 30410 207860 30480
rect 207640 30360 207860 30410
rect 204000 30350 208000 30360
rect 204000 30150 204020 30350
rect 204090 30150 204410 30350
rect 204480 30150 204520 30350
rect 204590 30150 204910 30350
rect 204980 30150 205020 30350
rect 205090 30150 205410 30350
rect 205480 30150 205520 30350
rect 205590 30150 205910 30350
rect 205980 30150 206020 30350
rect 206090 30150 206410 30350
rect 206480 30150 206520 30350
rect 206590 30150 206910 30350
rect 206980 30150 207020 30350
rect 207090 30150 207410 30350
rect 207480 30150 207520 30350
rect 207590 30150 207910 30350
rect 207980 30150 208000 30350
rect 204000 30140 208000 30150
rect 204140 30090 204360 30140
rect 204140 30020 204150 30090
rect 204350 30020 204360 30090
rect 204140 29980 204360 30020
rect 204140 29910 204150 29980
rect 204350 29910 204360 29980
rect 204140 29860 204360 29910
rect 204640 30090 204860 30140
rect 204640 30020 204650 30090
rect 204850 30020 204860 30090
rect 204640 29980 204860 30020
rect 204640 29910 204650 29980
rect 204850 29910 204860 29980
rect 204640 29860 204860 29910
rect 205140 30090 205360 30140
rect 205140 30020 205150 30090
rect 205350 30020 205360 30090
rect 205140 29980 205360 30020
rect 205140 29910 205150 29980
rect 205350 29910 205360 29980
rect 205140 29860 205360 29910
rect 205640 30090 205860 30140
rect 205640 30020 205650 30090
rect 205850 30020 205860 30090
rect 205640 29980 205860 30020
rect 205640 29910 205650 29980
rect 205850 29910 205860 29980
rect 205640 29860 205860 29910
rect 206140 30090 206360 30140
rect 206140 30020 206150 30090
rect 206350 30020 206360 30090
rect 206140 29980 206360 30020
rect 206140 29910 206150 29980
rect 206350 29910 206360 29980
rect 206140 29860 206360 29910
rect 206640 30090 206860 30140
rect 206640 30020 206650 30090
rect 206850 30020 206860 30090
rect 206640 29980 206860 30020
rect 206640 29910 206650 29980
rect 206850 29910 206860 29980
rect 206640 29860 206860 29910
rect 207140 30090 207360 30140
rect 207140 30020 207150 30090
rect 207350 30020 207360 30090
rect 207140 29980 207360 30020
rect 207140 29910 207150 29980
rect 207350 29910 207360 29980
rect 207140 29860 207360 29910
rect 207640 30090 207860 30140
rect 207640 30020 207650 30090
rect 207850 30020 207860 30090
rect 207640 29980 207860 30020
rect 207640 29910 207650 29980
rect 207850 29910 207860 29980
rect 207640 29860 207860 29910
rect 204000 29850 208000 29860
rect 204000 29650 204020 29850
rect 204090 29650 204410 29850
rect 204480 29650 204520 29850
rect 204590 29650 204910 29850
rect 204980 29650 205020 29850
rect 205090 29650 205410 29850
rect 205480 29650 205520 29850
rect 205590 29650 205910 29850
rect 205980 29650 206020 29850
rect 206090 29650 206410 29850
rect 206480 29650 206520 29850
rect 206590 29650 206910 29850
rect 206980 29650 207020 29850
rect 207090 29650 207410 29850
rect 207480 29650 207520 29850
rect 207590 29650 207910 29850
rect 207980 29650 208000 29850
rect 204000 29640 208000 29650
rect 204140 29590 204360 29640
rect 204140 29520 204150 29590
rect 204350 29520 204360 29590
rect 204140 29480 204360 29520
rect 204140 29410 204150 29480
rect 204350 29410 204360 29480
rect 204140 29360 204360 29410
rect 204640 29590 204860 29640
rect 204640 29520 204650 29590
rect 204850 29520 204860 29590
rect 204640 29480 204860 29520
rect 204640 29410 204650 29480
rect 204850 29410 204860 29480
rect 204640 29360 204860 29410
rect 205140 29590 205360 29640
rect 205140 29520 205150 29590
rect 205350 29520 205360 29590
rect 205140 29480 205360 29520
rect 205140 29410 205150 29480
rect 205350 29410 205360 29480
rect 205140 29360 205360 29410
rect 205640 29590 205860 29640
rect 205640 29520 205650 29590
rect 205850 29520 205860 29590
rect 205640 29480 205860 29520
rect 205640 29410 205650 29480
rect 205850 29410 205860 29480
rect 205640 29360 205860 29410
rect 206140 29590 206360 29640
rect 206140 29520 206150 29590
rect 206350 29520 206360 29590
rect 206140 29480 206360 29520
rect 206140 29410 206150 29480
rect 206350 29410 206360 29480
rect 206140 29360 206360 29410
rect 206640 29590 206860 29640
rect 206640 29520 206650 29590
rect 206850 29520 206860 29590
rect 206640 29480 206860 29520
rect 206640 29410 206650 29480
rect 206850 29410 206860 29480
rect 206640 29360 206860 29410
rect 207140 29590 207360 29640
rect 207140 29520 207150 29590
rect 207350 29520 207360 29590
rect 207140 29480 207360 29520
rect 207140 29410 207150 29480
rect 207350 29410 207360 29480
rect 207140 29360 207360 29410
rect 207640 29590 207860 29640
rect 207640 29520 207650 29590
rect 207850 29520 207860 29590
rect 207640 29480 207860 29520
rect 207640 29410 207650 29480
rect 207850 29410 207860 29480
rect 207640 29360 207860 29410
rect 204000 29350 208000 29360
rect 204000 29150 204020 29350
rect 204090 29150 204410 29350
rect 204480 29150 204520 29350
rect 204590 29150 204910 29350
rect 204980 29150 205020 29350
rect 205090 29150 205410 29350
rect 205480 29150 205520 29350
rect 205590 29150 205910 29350
rect 205980 29150 206020 29350
rect 206090 29150 206410 29350
rect 206480 29150 206520 29350
rect 206590 29150 206910 29350
rect 206980 29150 207020 29350
rect 207090 29150 207410 29350
rect 207480 29150 207520 29350
rect 207590 29150 207910 29350
rect 207980 29150 208000 29350
rect 204000 29140 208000 29150
rect 204140 29090 204360 29140
rect 204140 29020 204150 29090
rect 204350 29020 204360 29090
rect 204140 28980 204360 29020
rect 204140 28910 204150 28980
rect 204350 28910 204360 28980
rect 204140 28860 204360 28910
rect 204640 29090 204860 29140
rect 204640 29020 204650 29090
rect 204850 29020 204860 29090
rect 204640 28980 204860 29020
rect 204640 28910 204650 28980
rect 204850 28910 204860 28980
rect 204640 28860 204860 28910
rect 205140 29090 205360 29140
rect 205140 29020 205150 29090
rect 205350 29020 205360 29090
rect 205140 28980 205360 29020
rect 205140 28910 205150 28980
rect 205350 28910 205360 28980
rect 205140 28860 205360 28910
rect 205640 29090 205860 29140
rect 205640 29020 205650 29090
rect 205850 29020 205860 29090
rect 205640 28980 205860 29020
rect 205640 28910 205650 28980
rect 205850 28910 205860 28980
rect 205640 28860 205860 28910
rect 206140 29090 206360 29140
rect 206140 29020 206150 29090
rect 206350 29020 206360 29090
rect 206140 28980 206360 29020
rect 206140 28910 206150 28980
rect 206350 28910 206360 28980
rect 206140 28860 206360 28910
rect 206640 29090 206860 29140
rect 206640 29020 206650 29090
rect 206850 29020 206860 29090
rect 206640 28980 206860 29020
rect 206640 28910 206650 28980
rect 206850 28910 206860 28980
rect 206640 28860 206860 28910
rect 207140 29090 207360 29140
rect 207140 29020 207150 29090
rect 207350 29020 207360 29090
rect 207140 28980 207360 29020
rect 207140 28910 207150 28980
rect 207350 28910 207360 28980
rect 207140 28860 207360 28910
rect 207640 29090 207860 29140
rect 207640 29020 207650 29090
rect 207850 29020 207860 29090
rect 207640 28980 207860 29020
rect 207640 28910 207650 28980
rect 207850 28910 207860 28980
rect 207640 28860 207860 28910
rect 204000 28850 208000 28860
rect 204000 28650 204020 28850
rect 204090 28650 204410 28850
rect 204480 28650 204520 28850
rect 204590 28650 204910 28850
rect 204980 28650 205020 28850
rect 205090 28650 205410 28850
rect 205480 28650 205520 28850
rect 205590 28650 205910 28850
rect 205980 28650 206020 28850
rect 206090 28650 206410 28850
rect 206480 28650 206520 28850
rect 206590 28650 206910 28850
rect 206980 28650 207020 28850
rect 207090 28650 207410 28850
rect 207480 28650 207520 28850
rect 207590 28650 207910 28850
rect 207980 28650 208000 28850
rect 204000 28640 208000 28650
rect 204140 28590 204360 28640
rect 204140 28520 204150 28590
rect 204350 28520 204360 28590
rect 204140 28480 204360 28520
rect 204140 28410 204150 28480
rect 204350 28410 204360 28480
rect 204140 28360 204360 28410
rect 204640 28590 204860 28640
rect 204640 28520 204650 28590
rect 204850 28520 204860 28590
rect 204640 28480 204860 28520
rect 204640 28410 204650 28480
rect 204850 28410 204860 28480
rect 204640 28360 204860 28410
rect 205140 28590 205360 28640
rect 205140 28520 205150 28590
rect 205350 28520 205360 28590
rect 205140 28480 205360 28520
rect 205140 28410 205150 28480
rect 205350 28410 205360 28480
rect 205140 28360 205360 28410
rect 205640 28590 205860 28640
rect 205640 28520 205650 28590
rect 205850 28520 205860 28590
rect 205640 28480 205860 28520
rect 205640 28410 205650 28480
rect 205850 28410 205860 28480
rect 205640 28360 205860 28410
rect 206140 28590 206360 28640
rect 206140 28520 206150 28590
rect 206350 28520 206360 28590
rect 206140 28480 206360 28520
rect 206140 28410 206150 28480
rect 206350 28410 206360 28480
rect 206140 28360 206360 28410
rect 206640 28590 206860 28640
rect 206640 28520 206650 28590
rect 206850 28520 206860 28590
rect 206640 28480 206860 28520
rect 206640 28410 206650 28480
rect 206850 28410 206860 28480
rect 206640 28360 206860 28410
rect 207140 28590 207360 28640
rect 207140 28520 207150 28590
rect 207350 28520 207360 28590
rect 207140 28480 207360 28520
rect 207140 28410 207150 28480
rect 207350 28410 207360 28480
rect 207140 28360 207360 28410
rect 207640 28590 207860 28640
rect 207640 28520 207650 28590
rect 207850 28520 207860 28590
rect 207640 28480 207860 28520
rect 207640 28410 207650 28480
rect 207850 28410 207860 28480
rect 207640 28360 207860 28410
rect 204000 28350 208000 28360
rect 204000 28150 204020 28350
rect 204090 28150 204410 28350
rect 204480 28150 204520 28350
rect 204590 28150 204910 28350
rect 204980 28150 205020 28350
rect 205090 28150 205410 28350
rect 205480 28150 205520 28350
rect 205590 28150 205910 28350
rect 205980 28150 206020 28350
rect 206090 28150 206410 28350
rect 206480 28150 206520 28350
rect 206590 28150 206910 28350
rect 206980 28150 207020 28350
rect 207090 28150 207410 28350
rect 207480 28150 207520 28350
rect 207590 28150 207910 28350
rect 207980 28150 208000 28350
rect 204000 28140 208000 28150
rect 204140 28090 204360 28140
rect 204140 28020 204150 28090
rect 204350 28020 204360 28090
rect 204140 27980 204360 28020
rect 204140 27910 204150 27980
rect 204350 27910 204360 27980
rect 204140 27860 204360 27910
rect 204640 28090 204860 28140
rect 204640 28020 204650 28090
rect 204850 28020 204860 28090
rect 204640 27980 204860 28020
rect 204640 27910 204650 27980
rect 204850 27910 204860 27980
rect 204640 27860 204860 27910
rect 205140 28090 205360 28140
rect 205140 28020 205150 28090
rect 205350 28020 205360 28090
rect 205140 27980 205360 28020
rect 205140 27910 205150 27980
rect 205350 27910 205360 27980
rect 205140 27860 205360 27910
rect 205640 28090 205860 28140
rect 205640 28020 205650 28090
rect 205850 28020 205860 28090
rect 205640 27980 205860 28020
rect 205640 27910 205650 27980
rect 205850 27910 205860 27980
rect 205640 27860 205860 27910
rect 206140 28090 206360 28140
rect 206140 28020 206150 28090
rect 206350 28020 206360 28090
rect 206140 27980 206360 28020
rect 206140 27910 206150 27980
rect 206350 27910 206360 27980
rect 206140 27860 206360 27910
rect 206640 28090 206860 28140
rect 206640 28020 206650 28090
rect 206850 28020 206860 28090
rect 206640 27980 206860 28020
rect 206640 27910 206650 27980
rect 206850 27910 206860 27980
rect 206640 27860 206860 27910
rect 207140 28090 207360 28140
rect 207140 28020 207150 28090
rect 207350 28020 207360 28090
rect 207140 27980 207360 28020
rect 207140 27910 207150 27980
rect 207350 27910 207360 27980
rect 207140 27860 207360 27910
rect 207640 28090 207860 28140
rect 207640 28020 207650 28090
rect 207850 28020 207860 28090
rect 207640 27980 207860 28020
rect 207640 27910 207650 27980
rect 207850 27910 207860 27980
rect 207640 27860 207860 27910
rect 204000 27850 208000 27860
rect 204000 27650 204020 27850
rect 204090 27650 204410 27850
rect 204480 27650 204520 27850
rect 204590 27650 204910 27850
rect 204980 27650 205020 27850
rect 205090 27650 205410 27850
rect 205480 27650 205520 27850
rect 205590 27650 205910 27850
rect 205980 27650 206020 27850
rect 206090 27650 206410 27850
rect 206480 27650 206520 27850
rect 206590 27650 206910 27850
rect 206980 27650 207020 27850
rect 207090 27650 207410 27850
rect 207480 27650 207520 27850
rect 207590 27650 207910 27850
rect 207980 27650 208000 27850
rect 204000 27640 208000 27650
rect 204140 27590 204360 27640
rect 204140 27520 204150 27590
rect 204350 27520 204360 27590
rect 204140 27480 204360 27520
rect 204140 27410 204150 27480
rect 204350 27410 204360 27480
rect 204140 27360 204360 27410
rect 204640 27590 204860 27640
rect 204640 27520 204650 27590
rect 204850 27520 204860 27590
rect 204640 27480 204860 27520
rect 204640 27410 204650 27480
rect 204850 27410 204860 27480
rect 204640 27360 204860 27410
rect 205140 27590 205360 27640
rect 205140 27520 205150 27590
rect 205350 27520 205360 27590
rect 205140 27480 205360 27520
rect 205140 27410 205150 27480
rect 205350 27410 205360 27480
rect 205140 27360 205360 27410
rect 205640 27590 205860 27640
rect 205640 27520 205650 27590
rect 205850 27520 205860 27590
rect 205640 27480 205860 27520
rect 205640 27410 205650 27480
rect 205850 27410 205860 27480
rect 205640 27360 205860 27410
rect 206140 27590 206360 27640
rect 206140 27520 206150 27590
rect 206350 27520 206360 27590
rect 206140 27480 206360 27520
rect 206140 27410 206150 27480
rect 206350 27410 206360 27480
rect 206140 27360 206360 27410
rect 206640 27590 206860 27640
rect 206640 27520 206650 27590
rect 206850 27520 206860 27590
rect 206640 27480 206860 27520
rect 206640 27410 206650 27480
rect 206850 27410 206860 27480
rect 206640 27360 206860 27410
rect 207140 27590 207360 27640
rect 207140 27520 207150 27590
rect 207350 27520 207360 27590
rect 207140 27480 207360 27520
rect 207140 27410 207150 27480
rect 207350 27410 207360 27480
rect 207140 27360 207360 27410
rect 207640 27590 207860 27640
rect 207640 27520 207650 27590
rect 207850 27520 207860 27590
rect 207640 27480 207860 27520
rect 207640 27410 207650 27480
rect 207850 27410 207860 27480
rect 207640 27360 207860 27410
rect 204000 27350 208000 27360
rect 204000 27150 204020 27350
rect 204090 27150 204410 27350
rect 204480 27150 204520 27350
rect 204590 27150 204910 27350
rect 204980 27150 205020 27350
rect 205090 27150 205410 27350
rect 205480 27150 205520 27350
rect 205590 27150 205910 27350
rect 205980 27150 206020 27350
rect 206090 27150 206410 27350
rect 206480 27150 206520 27350
rect 206590 27150 206910 27350
rect 206980 27150 207020 27350
rect 207090 27150 207410 27350
rect 207480 27150 207520 27350
rect 207590 27150 207910 27350
rect 207980 27150 208000 27350
rect 204000 27140 208000 27150
rect 204140 27090 204360 27140
rect 204140 27020 204150 27090
rect 204350 27020 204360 27090
rect 204140 26980 204360 27020
rect 204140 26910 204150 26980
rect 204350 26910 204360 26980
rect 204140 26860 204360 26910
rect 204640 27090 204860 27140
rect 204640 27020 204650 27090
rect 204850 27020 204860 27090
rect 204640 26980 204860 27020
rect 204640 26910 204650 26980
rect 204850 26910 204860 26980
rect 204640 26860 204860 26910
rect 205140 27090 205360 27140
rect 205140 27020 205150 27090
rect 205350 27020 205360 27090
rect 205140 26980 205360 27020
rect 205140 26910 205150 26980
rect 205350 26910 205360 26980
rect 205140 26860 205360 26910
rect 205640 27090 205860 27140
rect 205640 27020 205650 27090
rect 205850 27020 205860 27090
rect 205640 26980 205860 27020
rect 205640 26910 205650 26980
rect 205850 26910 205860 26980
rect 205640 26860 205860 26910
rect 206140 27090 206360 27140
rect 206140 27020 206150 27090
rect 206350 27020 206360 27090
rect 206140 26980 206360 27020
rect 206140 26910 206150 26980
rect 206350 26910 206360 26980
rect 206140 26860 206360 26910
rect 206640 27090 206860 27140
rect 206640 27020 206650 27090
rect 206850 27020 206860 27090
rect 206640 26980 206860 27020
rect 206640 26910 206650 26980
rect 206850 26910 206860 26980
rect 206640 26860 206860 26910
rect 207140 27090 207360 27140
rect 207140 27020 207150 27090
rect 207350 27020 207360 27090
rect 207140 26980 207360 27020
rect 207140 26910 207150 26980
rect 207350 26910 207360 26980
rect 207140 26860 207360 26910
rect 207640 27090 207860 27140
rect 207640 27020 207650 27090
rect 207850 27020 207860 27090
rect 207640 26980 207860 27020
rect 207640 26910 207650 26980
rect 207850 26910 207860 26980
rect 207640 26860 207860 26910
rect 204000 26850 208000 26860
rect 204000 26650 204020 26850
rect 204090 26650 204410 26850
rect 204480 26650 204520 26850
rect 204590 26650 204910 26850
rect 204980 26650 205020 26850
rect 205090 26650 205410 26850
rect 205480 26650 205520 26850
rect 205590 26650 205910 26850
rect 205980 26650 206020 26850
rect 206090 26650 206410 26850
rect 206480 26650 206520 26850
rect 206590 26650 206910 26850
rect 206980 26650 207020 26850
rect 207090 26650 207410 26850
rect 207480 26650 207520 26850
rect 207590 26650 207910 26850
rect 207980 26650 208000 26850
rect 204000 26640 208000 26650
rect 204140 26590 204360 26640
rect 204140 26520 204150 26590
rect 204350 26520 204360 26590
rect 204140 26480 204360 26520
rect 204140 26410 204150 26480
rect 204350 26410 204360 26480
rect 204140 26360 204360 26410
rect 204640 26590 204860 26640
rect 204640 26520 204650 26590
rect 204850 26520 204860 26590
rect 204640 26480 204860 26520
rect 204640 26410 204650 26480
rect 204850 26410 204860 26480
rect 204640 26360 204860 26410
rect 205140 26590 205360 26640
rect 205140 26520 205150 26590
rect 205350 26520 205360 26590
rect 205140 26480 205360 26520
rect 205140 26410 205150 26480
rect 205350 26410 205360 26480
rect 205140 26360 205360 26410
rect 205640 26590 205860 26640
rect 205640 26520 205650 26590
rect 205850 26520 205860 26590
rect 205640 26480 205860 26520
rect 205640 26410 205650 26480
rect 205850 26410 205860 26480
rect 205640 26360 205860 26410
rect 206140 26590 206360 26640
rect 206140 26520 206150 26590
rect 206350 26520 206360 26590
rect 206140 26480 206360 26520
rect 206140 26410 206150 26480
rect 206350 26410 206360 26480
rect 206140 26360 206360 26410
rect 206640 26590 206860 26640
rect 206640 26520 206650 26590
rect 206850 26520 206860 26590
rect 206640 26480 206860 26520
rect 206640 26410 206650 26480
rect 206850 26410 206860 26480
rect 206640 26360 206860 26410
rect 207140 26590 207360 26640
rect 207140 26520 207150 26590
rect 207350 26520 207360 26590
rect 207140 26480 207360 26520
rect 207140 26410 207150 26480
rect 207350 26410 207360 26480
rect 207140 26360 207360 26410
rect 207640 26590 207860 26640
rect 207640 26520 207650 26590
rect 207850 26520 207860 26590
rect 207640 26480 207860 26520
rect 207640 26410 207650 26480
rect 207850 26410 207860 26480
rect 207640 26360 207860 26410
rect 204000 26350 208000 26360
rect 204000 26150 204020 26350
rect 204090 26150 204410 26350
rect 204480 26150 204520 26350
rect 204590 26150 204910 26350
rect 204980 26150 205020 26350
rect 205090 26150 205410 26350
rect 205480 26150 205520 26350
rect 205590 26150 205910 26350
rect 205980 26150 206020 26350
rect 206090 26150 206410 26350
rect 206480 26150 206520 26350
rect 206590 26150 206910 26350
rect 206980 26150 207020 26350
rect 207090 26150 207410 26350
rect 207480 26150 207520 26350
rect 207590 26150 207910 26350
rect 207980 26150 208000 26350
rect 204000 26140 208000 26150
rect 204140 26090 204360 26140
rect 204140 26020 204150 26090
rect 204350 26020 204360 26090
rect 204140 25980 204360 26020
rect 204140 25910 204150 25980
rect 204350 25910 204360 25980
rect 204140 25860 204360 25910
rect 204640 26090 204860 26140
rect 204640 26020 204650 26090
rect 204850 26020 204860 26090
rect 204640 25980 204860 26020
rect 204640 25910 204650 25980
rect 204850 25910 204860 25980
rect 204640 25860 204860 25910
rect 205140 26090 205360 26140
rect 205140 26020 205150 26090
rect 205350 26020 205360 26090
rect 205140 25980 205360 26020
rect 205140 25910 205150 25980
rect 205350 25910 205360 25980
rect 205140 25860 205360 25910
rect 205640 26090 205860 26140
rect 205640 26020 205650 26090
rect 205850 26020 205860 26090
rect 205640 25980 205860 26020
rect 205640 25910 205650 25980
rect 205850 25910 205860 25980
rect 205640 25860 205860 25910
rect 206140 26090 206360 26140
rect 206140 26020 206150 26090
rect 206350 26020 206360 26090
rect 206140 25980 206360 26020
rect 206140 25910 206150 25980
rect 206350 25910 206360 25980
rect 206140 25860 206360 25910
rect 206640 26090 206860 26140
rect 206640 26020 206650 26090
rect 206850 26020 206860 26090
rect 206640 25980 206860 26020
rect 206640 25910 206650 25980
rect 206850 25910 206860 25980
rect 206640 25860 206860 25910
rect 207140 26090 207360 26140
rect 207140 26020 207150 26090
rect 207350 26020 207360 26090
rect 207140 25980 207360 26020
rect 207140 25910 207150 25980
rect 207350 25910 207360 25980
rect 207140 25860 207360 25910
rect 207640 26090 207860 26140
rect 207640 26020 207650 26090
rect 207850 26020 207860 26090
rect 207640 25980 207860 26020
rect 207640 25910 207650 25980
rect 207850 25910 207860 25980
rect 207640 25860 207860 25910
rect 204000 25850 208000 25860
rect 204000 25650 204020 25850
rect 204090 25650 204410 25850
rect 204480 25650 204520 25850
rect 204590 25650 204910 25850
rect 204980 25650 205020 25850
rect 205090 25650 205410 25850
rect 205480 25650 205520 25850
rect 205590 25650 205910 25850
rect 205980 25650 206020 25850
rect 206090 25650 206410 25850
rect 206480 25650 206520 25850
rect 206590 25650 206910 25850
rect 206980 25650 207020 25850
rect 207090 25650 207410 25850
rect 207480 25650 207520 25850
rect 207590 25650 207910 25850
rect 207980 25650 208000 25850
rect 204000 25640 208000 25650
rect 204140 25590 204360 25640
rect 204140 25520 204150 25590
rect 204350 25520 204360 25590
rect 204140 25480 204360 25520
rect 204140 25410 204150 25480
rect 204350 25410 204360 25480
rect 204140 25360 204360 25410
rect 204640 25590 204860 25640
rect 204640 25520 204650 25590
rect 204850 25520 204860 25590
rect 204640 25480 204860 25520
rect 204640 25410 204650 25480
rect 204850 25410 204860 25480
rect 204640 25360 204860 25410
rect 205140 25590 205360 25640
rect 205140 25520 205150 25590
rect 205350 25520 205360 25590
rect 205140 25480 205360 25520
rect 205140 25410 205150 25480
rect 205350 25410 205360 25480
rect 205140 25360 205360 25410
rect 205640 25590 205860 25640
rect 205640 25520 205650 25590
rect 205850 25520 205860 25590
rect 205640 25480 205860 25520
rect 205640 25410 205650 25480
rect 205850 25410 205860 25480
rect 205640 25360 205860 25410
rect 206140 25590 206360 25640
rect 206140 25520 206150 25590
rect 206350 25520 206360 25590
rect 206140 25480 206360 25520
rect 206140 25410 206150 25480
rect 206350 25410 206360 25480
rect 206140 25360 206360 25410
rect 206640 25590 206860 25640
rect 206640 25520 206650 25590
rect 206850 25520 206860 25590
rect 206640 25480 206860 25520
rect 206640 25410 206650 25480
rect 206850 25410 206860 25480
rect 206640 25360 206860 25410
rect 207140 25590 207360 25640
rect 207140 25520 207150 25590
rect 207350 25520 207360 25590
rect 207140 25480 207360 25520
rect 207140 25410 207150 25480
rect 207350 25410 207360 25480
rect 207140 25360 207360 25410
rect 207640 25590 207860 25640
rect 207640 25520 207650 25590
rect 207850 25520 207860 25590
rect 207640 25480 207860 25520
rect 207640 25410 207650 25480
rect 207850 25410 207860 25480
rect 207640 25360 207860 25410
rect 204000 25350 208000 25360
rect 204000 25150 204020 25350
rect 204090 25150 204410 25350
rect 204480 25150 204520 25350
rect 204590 25150 204910 25350
rect 204980 25150 205020 25350
rect 205090 25150 205410 25350
rect 205480 25150 205520 25350
rect 205590 25150 205910 25350
rect 205980 25150 206020 25350
rect 206090 25150 206410 25350
rect 206480 25150 206520 25350
rect 206590 25150 206910 25350
rect 206980 25150 207020 25350
rect 207090 25150 207410 25350
rect 207480 25150 207520 25350
rect 207590 25150 207910 25350
rect 207980 25150 208000 25350
rect 204000 25140 208000 25150
rect 204140 25090 204360 25140
rect 204140 25020 204150 25090
rect 204350 25020 204360 25090
rect 204140 24980 204360 25020
rect 204140 24910 204150 24980
rect 204350 24910 204360 24980
rect 204140 24860 204360 24910
rect 204640 25090 204860 25140
rect 204640 25020 204650 25090
rect 204850 25020 204860 25090
rect 204640 24980 204860 25020
rect 204640 24910 204650 24980
rect 204850 24910 204860 24980
rect 204640 24860 204860 24910
rect 205140 25090 205360 25140
rect 205140 25020 205150 25090
rect 205350 25020 205360 25090
rect 205140 24980 205360 25020
rect 205140 24910 205150 24980
rect 205350 24910 205360 24980
rect 205140 24860 205360 24910
rect 205640 25090 205860 25140
rect 205640 25020 205650 25090
rect 205850 25020 205860 25090
rect 205640 24980 205860 25020
rect 205640 24910 205650 24980
rect 205850 24910 205860 24980
rect 205640 24860 205860 24910
rect 206140 25090 206360 25140
rect 206140 25020 206150 25090
rect 206350 25020 206360 25090
rect 206140 24980 206360 25020
rect 206140 24910 206150 24980
rect 206350 24910 206360 24980
rect 206140 24860 206360 24910
rect 206640 25090 206860 25140
rect 206640 25020 206650 25090
rect 206850 25020 206860 25090
rect 206640 24980 206860 25020
rect 206640 24910 206650 24980
rect 206850 24910 206860 24980
rect 206640 24860 206860 24910
rect 207140 25090 207360 25140
rect 207140 25020 207150 25090
rect 207350 25020 207360 25090
rect 207140 24980 207360 25020
rect 207140 24910 207150 24980
rect 207350 24910 207360 24980
rect 207140 24860 207360 24910
rect 207640 25090 207860 25140
rect 207640 25020 207650 25090
rect 207850 25020 207860 25090
rect 207640 24980 207860 25020
rect 207640 24910 207650 24980
rect 207850 24910 207860 24980
rect 207640 24860 207860 24910
rect 204000 24850 208000 24860
rect 204000 24650 204020 24850
rect 204090 24650 204410 24850
rect 204480 24650 204520 24850
rect 204590 24650 204910 24850
rect 204980 24650 205020 24850
rect 205090 24650 205410 24850
rect 205480 24650 205520 24850
rect 205590 24650 205910 24850
rect 205980 24650 206020 24850
rect 206090 24650 206410 24850
rect 206480 24650 206520 24850
rect 206590 24650 206910 24850
rect 206980 24650 207020 24850
rect 207090 24650 207410 24850
rect 207480 24650 207520 24850
rect 207590 24650 207910 24850
rect 207980 24650 208000 24850
rect 204000 24640 208000 24650
rect 204140 24590 204360 24640
rect 204140 24520 204150 24590
rect 204350 24520 204360 24590
rect 204140 24480 204360 24520
rect 204140 24410 204150 24480
rect 204350 24410 204360 24480
rect 204140 24360 204360 24410
rect 204640 24590 204860 24640
rect 204640 24520 204650 24590
rect 204850 24520 204860 24590
rect 204640 24480 204860 24520
rect 204640 24410 204650 24480
rect 204850 24410 204860 24480
rect 204640 24360 204860 24410
rect 205140 24590 205360 24640
rect 205140 24520 205150 24590
rect 205350 24520 205360 24590
rect 205140 24480 205360 24520
rect 205140 24410 205150 24480
rect 205350 24410 205360 24480
rect 205140 24360 205360 24410
rect 205640 24590 205860 24640
rect 205640 24520 205650 24590
rect 205850 24520 205860 24590
rect 205640 24480 205860 24520
rect 205640 24410 205650 24480
rect 205850 24410 205860 24480
rect 205640 24360 205860 24410
rect 206140 24590 206360 24640
rect 206140 24520 206150 24590
rect 206350 24520 206360 24590
rect 206140 24480 206360 24520
rect 206140 24410 206150 24480
rect 206350 24410 206360 24480
rect 206140 24360 206360 24410
rect 206640 24590 206860 24640
rect 206640 24520 206650 24590
rect 206850 24520 206860 24590
rect 206640 24480 206860 24520
rect 206640 24410 206650 24480
rect 206850 24410 206860 24480
rect 206640 24360 206860 24410
rect 207140 24590 207360 24640
rect 207140 24520 207150 24590
rect 207350 24520 207360 24590
rect 207140 24480 207360 24520
rect 207140 24410 207150 24480
rect 207350 24410 207360 24480
rect 207140 24360 207360 24410
rect 207640 24590 207860 24640
rect 207640 24520 207650 24590
rect 207850 24520 207860 24590
rect 207640 24480 207860 24520
rect 207640 24410 207650 24480
rect 207850 24410 207860 24480
rect 207640 24360 207860 24410
rect 204000 24350 208000 24360
rect 204000 24150 204020 24350
rect 204090 24150 204410 24350
rect 204480 24150 204520 24350
rect 204590 24150 204910 24350
rect 204980 24150 205020 24350
rect 205090 24150 205410 24350
rect 205480 24150 205520 24350
rect 205590 24150 205910 24350
rect 205980 24150 206020 24350
rect 206090 24150 206410 24350
rect 206480 24150 206520 24350
rect 206590 24150 206910 24350
rect 206980 24150 207020 24350
rect 207090 24150 207410 24350
rect 207480 24150 207520 24350
rect 207590 24150 207910 24350
rect 207980 24150 208000 24350
rect 204000 24140 208000 24150
rect 204140 24090 204360 24140
rect 204140 24020 204150 24090
rect 204350 24020 204360 24090
rect 204140 23980 204360 24020
rect 204140 23910 204150 23980
rect 204350 23910 204360 23980
rect 204140 23860 204360 23910
rect 204640 24090 204860 24140
rect 204640 24020 204650 24090
rect 204850 24020 204860 24090
rect 204640 23980 204860 24020
rect 204640 23910 204650 23980
rect 204850 23910 204860 23980
rect 204640 23860 204860 23910
rect 205140 24090 205360 24140
rect 205140 24020 205150 24090
rect 205350 24020 205360 24090
rect 205140 23980 205360 24020
rect 205140 23910 205150 23980
rect 205350 23910 205360 23980
rect 205140 23860 205360 23910
rect 205640 24090 205860 24140
rect 205640 24020 205650 24090
rect 205850 24020 205860 24090
rect 205640 23980 205860 24020
rect 205640 23910 205650 23980
rect 205850 23910 205860 23980
rect 205640 23860 205860 23910
rect 206140 24090 206360 24140
rect 206140 24020 206150 24090
rect 206350 24020 206360 24090
rect 206140 23980 206360 24020
rect 206140 23910 206150 23980
rect 206350 23910 206360 23980
rect 206140 23860 206360 23910
rect 206640 24090 206860 24140
rect 206640 24020 206650 24090
rect 206850 24020 206860 24090
rect 206640 23980 206860 24020
rect 206640 23910 206650 23980
rect 206850 23910 206860 23980
rect 206640 23860 206860 23910
rect 207140 24090 207360 24140
rect 207140 24020 207150 24090
rect 207350 24020 207360 24090
rect 207140 23980 207360 24020
rect 207140 23910 207150 23980
rect 207350 23910 207360 23980
rect 207140 23860 207360 23910
rect 207640 24090 207860 24140
rect 207640 24020 207650 24090
rect 207850 24020 207860 24090
rect 207640 23980 207860 24020
rect 207640 23910 207650 23980
rect 207850 23910 207860 23980
rect 207640 23860 207860 23910
rect 204000 23850 208000 23860
rect 204000 23650 204020 23850
rect 204090 23650 204410 23850
rect 204480 23650 204520 23850
rect 204590 23650 204910 23850
rect 204980 23650 205020 23850
rect 205090 23650 205410 23850
rect 205480 23650 205520 23850
rect 205590 23650 205910 23850
rect 205980 23650 206020 23850
rect 206090 23650 206410 23850
rect 206480 23650 206520 23850
rect 206590 23650 206910 23850
rect 206980 23650 207020 23850
rect 207090 23650 207410 23850
rect 207480 23650 207520 23850
rect 207590 23650 207910 23850
rect 207980 23650 208000 23850
rect 204000 23640 208000 23650
rect 204140 23590 204360 23640
rect 204140 23520 204150 23590
rect 204350 23520 204360 23590
rect 204140 23480 204360 23520
rect 204140 23410 204150 23480
rect 204350 23410 204360 23480
rect 204140 23360 204360 23410
rect 204640 23590 204860 23640
rect 204640 23520 204650 23590
rect 204850 23520 204860 23590
rect 204640 23480 204860 23520
rect 204640 23410 204650 23480
rect 204850 23410 204860 23480
rect 204640 23360 204860 23410
rect 205140 23590 205360 23640
rect 205140 23520 205150 23590
rect 205350 23520 205360 23590
rect 205140 23480 205360 23520
rect 205140 23410 205150 23480
rect 205350 23410 205360 23480
rect 205140 23360 205360 23410
rect 205640 23590 205860 23640
rect 205640 23520 205650 23590
rect 205850 23520 205860 23590
rect 205640 23480 205860 23520
rect 205640 23410 205650 23480
rect 205850 23410 205860 23480
rect 205640 23360 205860 23410
rect 206140 23590 206360 23640
rect 206140 23520 206150 23590
rect 206350 23520 206360 23590
rect 206140 23480 206360 23520
rect 206140 23410 206150 23480
rect 206350 23410 206360 23480
rect 206140 23360 206360 23410
rect 206640 23590 206860 23640
rect 206640 23520 206650 23590
rect 206850 23520 206860 23590
rect 206640 23480 206860 23520
rect 206640 23410 206650 23480
rect 206850 23410 206860 23480
rect 206640 23360 206860 23410
rect 207140 23590 207360 23640
rect 207140 23520 207150 23590
rect 207350 23520 207360 23590
rect 207140 23480 207360 23520
rect 207140 23410 207150 23480
rect 207350 23410 207360 23480
rect 207140 23360 207360 23410
rect 207640 23590 207860 23640
rect 207640 23520 207650 23590
rect 207850 23520 207860 23590
rect 207640 23480 207860 23520
rect 207640 23410 207650 23480
rect 207850 23410 207860 23480
rect 207640 23360 207860 23410
rect 204000 23350 208000 23360
rect 204000 23150 204020 23350
rect 204090 23150 204410 23350
rect 204480 23150 204520 23350
rect 204590 23150 204910 23350
rect 204980 23150 205020 23350
rect 205090 23150 205410 23350
rect 205480 23150 205520 23350
rect 205590 23150 205910 23350
rect 205980 23150 206020 23350
rect 206090 23150 206410 23350
rect 206480 23150 206520 23350
rect 206590 23150 206910 23350
rect 206980 23150 207020 23350
rect 207090 23150 207410 23350
rect 207480 23150 207520 23350
rect 207590 23150 207910 23350
rect 207980 23150 208000 23350
rect 204000 23140 208000 23150
rect 204140 23090 204360 23140
rect 204140 23020 204150 23090
rect 204350 23020 204360 23090
rect 204140 22980 204360 23020
rect 204140 22910 204150 22980
rect 204350 22910 204360 22980
rect 204140 22860 204360 22910
rect 204640 23090 204860 23140
rect 204640 23020 204650 23090
rect 204850 23020 204860 23090
rect 204640 22980 204860 23020
rect 204640 22910 204650 22980
rect 204850 22910 204860 22980
rect 204640 22860 204860 22910
rect 205140 23090 205360 23140
rect 205140 23020 205150 23090
rect 205350 23020 205360 23090
rect 205140 22980 205360 23020
rect 205140 22910 205150 22980
rect 205350 22910 205360 22980
rect 205140 22860 205360 22910
rect 205640 23090 205860 23140
rect 205640 23020 205650 23090
rect 205850 23020 205860 23090
rect 205640 22980 205860 23020
rect 205640 22910 205650 22980
rect 205850 22910 205860 22980
rect 205640 22860 205860 22910
rect 206140 23090 206360 23140
rect 206140 23020 206150 23090
rect 206350 23020 206360 23090
rect 206140 22980 206360 23020
rect 206140 22910 206150 22980
rect 206350 22910 206360 22980
rect 206140 22860 206360 22910
rect 206640 23090 206860 23140
rect 206640 23020 206650 23090
rect 206850 23020 206860 23090
rect 206640 22980 206860 23020
rect 206640 22910 206650 22980
rect 206850 22910 206860 22980
rect 206640 22860 206860 22910
rect 207140 23090 207360 23140
rect 207140 23020 207150 23090
rect 207350 23020 207360 23090
rect 207140 22980 207360 23020
rect 207140 22910 207150 22980
rect 207350 22910 207360 22980
rect 207140 22860 207360 22910
rect 207640 23090 207860 23140
rect 207640 23020 207650 23090
rect 207850 23020 207860 23090
rect 207640 22980 207860 23020
rect 207640 22910 207650 22980
rect 207850 22910 207860 22980
rect 207640 22860 207860 22910
rect 204000 22850 208000 22860
rect 204000 22650 204020 22850
rect 204090 22650 204410 22850
rect 204480 22650 204520 22850
rect 204590 22650 204910 22850
rect 204980 22650 205020 22850
rect 205090 22650 205410 22850
rect 205480 22650 205520 22850
rect 205590 22650 205910 22850
rect 205980 22650 206020 22850
rect 206090 22650 206410 22850
rect 206480 22650 206520 22850
rect 206590 22650 206910 22850
rect 206980 22650 207020 22850
rect 207090 22650 207410 22850
rect 207480 22650 207520 22850
rect 207590 22650 207910 22850
rect 207980 22650 208000 22850
rect 204000 22640 208000 22650
rect 204140 22590 204360 22640
rect 204140 22520 204150 22590
rect 204350 22520 204360 22590
rect 204140 22480 204360 22520
rect 204140 22410 204150 22480
rect 204350 22410 204360 22480
rect 204140 22360 204360 22410
rect 204640 22590 204860 22640
rect 204640 22520 204650 22590
rect 204850 22520 204860 22590
rect 204640 22480 204860 22520
rect 204640 22410 204650 22480
rect 204850 22410 204860 22480
rect 204640 22360 204860 22410
rect 205140 22590 205360 22640
rect 205140 22520 205150 22590
rect 205350 22520 205360 22590
rect 205140 22480 205360 22520
rect 205140 22410 205150 22480
rect 205350 22410 205360 22480
rect 205140 22360 205360 22410
rect 205640 22590 205860 22640
rect 205640 22520 205650 22590
rect 205850 22520 205860 22590
rect 205640 22480 205860 22520
rect 205640 22410 205650 22480
rect 205850 22410 205860 22480
rect 205640 22360 205860 22410
rect 206140 22590 206360 22640
rect 206140 22520 206150 22590
rect 206350 22520 206360 22590
rect 206140 22480 206360 22520
rect 206140 22410 206150 22480
rect 206350 22410 206360 22480
rect 206140 22360 206360 22410
rect 206640 22590 206860 22640
rect 206640 22520 206650 22590
rect 206850 22520 206860 22590
rect 206640 22480 206860 22520
rect 206640 22410 206650 22480
rect 206850 22410 206860 22480
rect 206640 22360 206860 22410
rect 207140 22590 207360 22640
rect 207140 22520 207150 22590
rect 207350 22520 207360 22590
rect 207140 22480 207360 22520
rect 207140 22410 207150 22480
rect 207350 22410 207360 22480
rect 207140 22360 207360 22410
rect 207640 22590 207860 22640
rect 207640 22520 207650 22590
rect 207850 22520 207860 22590
rect 207640 22480 207860 22520
rect 207640 22410 207650 22480
rect 207850 22410 207860 22480
rect 207640 22360 207860 22410
rect 204000 22350 208000 22360
rect 204000 22150 204020 22350
rect 204090 22150 204410 22350
rect 204480 22150 204520 22350
rect 204590 22150 204910 22350
rect 204980 22150 205020 22350
rect 205090 22150 205410 22350
rect 205480 22150 205520 22350
rect 205590 22150 205910 22350
rect 205980 22150 206020 22350
rect 206090 22150 206410 22350
rect 206480 22150 206520 22350
rect 206590 22150 206910 22350
rect 206980 22150 207020 22350
rect 207090 22150 207410 22350
rect 207480 22150 207520 22350
rect 207590 22150 207910 22350
rect 207980 22150 208000 22350
rect 204000 22140 208000 22150
rect 204140 22090 204360 22140
rect 204140 22020 204150 22090
rect 204350 22020 204360 22090
rect 204140 21980 204360 22020
rect 204140 21910 204150 21980
rect 204350 21910 204360 21980
rect 204140 21860 204360 21910
rect 204640 22090 204860 22140
rect 204640 22020 204650 22090
rect 204850 22020 204860 22090
rect 204640 21980 204860 22020
rect 204640 21910 204650 21980
rect 204850 21910 204860 21980
rect 204640 21860 204860 21910
rect 205140 22090 205360 22140
rect 205140 22020 205150 22090
rect 205350 22020 205360 22090
rect 205140 21980 205360 22020
rect 205140 21910 205150 21980
rect 205350 21910 205360 21980
rect 205140 21860 205360 21910
rect 205640 22090 205860 22140
rect 205640 22020 205650 22090
rect 205850 22020 205860 22090
rect 205640 21980 205860 22020
rect 205640 21910 205650 21980
rect 205850 21910 205860 21980
rect 205640 21860 205860 21910
rect 206140 22090 206360 22140
rect 206140 22020 206150 22090
rect 206350 22020 206360 22090
rect 206140 21980 206360 22020
rect 206140 21910 206150 21980
rect 206350 21910 206360 21980
rect 206140 21860 206360 21910
rect 206640 22090 206860 22140
rect 206640 22020 206650 22090
rect 206850 22020 206860 22090
rect 206640 21980 206860 22020
rect 206640 21910 206650 21980
rect 206850 21910 206860 21980
rect 206640 21860 206860 21910
rect 207140 22090 207360 22140
rect 207140 22020 207150 22090
rect 207350 22020 207360 22090
rect 207140 21980 207360 22020
rect 207140 21910 207150 21980
rect 207350 21910 207360 21980
rect 207140 21860 207360 21910
rect 207640 22090 207860 22140
rect 207640 22020 207650 22090
rect 207850 22020 207860 22090
rect 207640 21980 207860 22020
rect 207640 21910 207650 21980
rect 207850 21910 207860 21980
rect 207640 21860 207860 21910
rect 204000 21850 208000 21860
rect 204000 21650 204020 21850
rect 204090 21650 204410 21850
rect 204480 21650 204520 21850
rect 204590 21650 204910 21850
rect 204980 21650 205020 21850
rect 205090 21650 205410 21850
rect 205480 21650 205520 21850
rect 205590 21650 205910 21850
rect 205980 21650 206020 21850
rect 206090 21650 206410 21850
rect 206480 21650 206520 21850
rect 206590 21650 206910 21850
rect 206980 21650 207020 21850
rect 207090 21650 207410 21850
rect 207480 21650 207520 21850
rect 207590 21650 207910 21850
rect 207980 21650 208000 21850
rect 204000 21640 208000 21650
rect 204140 21590 204360 21640
rect 204140 21520 204150 21590
rect 204350 21520 204360 21590
rect 204140 21480 204360 21520
rect 204140 21410 204150 21480
rect 204350 21410 204360 21480
rect 204140 21360 204360 21410
rect 204640 21590 204860 21640
rect 204640 21520 204650 21590
rect 204850 21520 204860 21590
rect 204640 21480 204860 21520
rect 204640 21410 204650 21480
rect 204850 21410 204860 21480
rect 204640 21360 204860 21410
rect 205140 21590 205360 21640
rect 205140 21520 205150 21590
rect 205350 21520 205360 21590
rect 205140 21480 205360 21520
rect 205140 21410 205150 21480
rect 205350 21410 205360 21480
rect 205140 21360 205360 21410
rect 205640 21590 205860 21640
rect 205640 21520 205650 21590
rect 205850 21520 205860 21590
rect 205640 21480 205860 21520
rect 205640 21410 205650 21480
rect 205850 21410 205860 21480
rect 205640 21360 205860 21410
rect 206140 21590 206360 21640
rect 206140 21520 206150 21590
rect 206350 21520 206360 21590
rect 206140 21480 206360 21520
rect 206140 21410 206150 21480
rect 206350 21410 206360 21480
rect 206140 21360 206360 21410
rect 206640 21590 206860 21640
rect 206640 21520 206650 21590
rect 206850 21520 206860 21590
rect 206640 21480 206860 21520
rect 206640 21410 206650 21480
rect 206850 21410 206860 21480
rect 206640 21360 206860 21410
rect 207140 21590 207360 21640
rect 207140 21520 207150 21590
rect 207350 21520 207360 21590
rect 207140 21480 207360 21520
rect 207140 21410 207150 21480
rect 207350 21410 207360 21480
rect 207140 21360 207360 21410
rect 207640 21590 207860 21640
rect 207640 21520 207650 21590
rect 207850 21520 207860 21590
rect 207640 21480 207860 21520
rect 207640 21410 207650 21480
rect 207850 21410 207860 21480
rect 207640 21360 207860 21410
rect 204000 21350 208000 21360
rect 204000 21150 204020 21350
rect 204090 21150 204410 21350
rect 204480 21150 204520 21350
rect 204590 21150 204910 21350
rect 204980 21150 205020 21350
rect 205090 21150 205410 21350
rect 205480 21150 205520 21350
rect 205590 21150 205910 21350
rect 205980 21150 206020 21350
rect 206090 21150 206410 21350
rect 206480 21150 206520 21350
rect 206590 21150 206910 21350
rect 206980 21150 207020 21350
rect 207090 21150 207410 21350
rect 207480 21150 207520 21350
rect 207590 21150 207910 21350
rect 207980 21150 208000 21350
rect 204000 21140 208000 21150
rect 204140 21090 204360 21140
rect 204140 21020 204150 21090
rect 204350 21020 204360 21090
rect 204140 20980 204360 21020
rect 204140 20910 204150 20980
rect 204350 20910 204360 20980
rect 204140 20860 204360 20910
rect 204640 21090 204860 21140
rect 204640 21020 204650 21090
rect 204850 21020 204860 21090
rect 204640 20980 204860 21020
rect 204640 20910 204650 20980
rect 204850 20910 204860 20980
rect 204640 20860 204860 20910
rect 205140 21090 205360 21140
rect 205140 21020 205150 21090
rect 205350 21020 205360 21090
rect 205140 20980 205360 21020
rect 205140 20910 205150 20980
rect 205350 20910 205360 20980
rect 205140 20860 205360 20910
rect 205640 21090 205860 21140
rect 205640 21020 205650 21090
rect 205850 21020 205860 21090
rect 205640 20980 205860 21020
rect 205640 20910 205650 20980
rect 205850 20910 205860 20980
rect 205640 20860 205860 20910
rect 206140 21090 206360 21140
rect 206140 21020 206150 21090
rect 206350 21020 206360 21090
rect 206140 20980 206360 21020
rect 206140 20910 206150 20980
rect 206350 20910 206360 20980
rect 206140 20860 206360 20910
rect 206640 21090 206860 21140
rect 206640 21020 206650 21090
rect 206850 21020 206860 21090
rect 206640 20980 206860 21020
rect 206640 20910 206650 20980
rect 206850 20910 206860 20980
rect 206640 20860 206860 20910
rect 207140 21090 207360 21140
rect 207140 21020 207150 21090
rect 207350 21020 207360 21090
rect 207140 20980 207360 21020
rect 207140 20910 207150 20980
rect 207350 20910 207360 20980
rect 207140 20860 207360 20910
rect 207640 21090 207860 21140
rect 207640 21020 207650 21090
rect 207850 21020 207860 21090
rect 207640 20980 207860 21020
rect 207640 20910 207650 20980
rect 207850 20910 207860 20980
rect 207640 20860 207860 20910
rect 204000 20850 208000 20860
rect 204000 20650 204020 20850
rect 204090 20650 204410 20850
rect 204480 20650 204520 20850
rect 204590 20650 204910 20850
rect 204980 20650 205020 20850
rect 205090 20650 205410 20850
rect 205480 20650 205520 20850
rect 205590 20650 205910 20850
rect 205980 20650 206020 20850
rect 206090 20650 206410 20850
rect 206480 20650 206520 20850
rect 206590 20650 206910 20850
rect 206980 20650 207020 20850
rect 207090 20650 207410 20850
rect 207480 20650 207520 20850
rect 207590 20650 207910 20850
rect 207980 20650 208000 20850
rect 204000 20640 208000 20650
rect 204140 20590 204360 20640
rect 204140 20520 204150 20590
rect 204350 20520 204360 20590
rect 204140 20480 204360 20520
rect 204140 20410 204150 20480
rect 204350 20410 204360 20480
rect 204140 20360 204360 20410
rect 204640 20590 204860 20640
rect 204640 20520 204650 20590
rect 204850 20520 204860 20590
rect 204640 20480 204860 20520
rect 204640 20410 204650 20480
rect 204850 20410 204860 20480
rect 204640 20360 204860 20410
rect 205140 20590 205360 20640
rect 205140 20520 205150 20590
rect 205350 20520 205360 20590
rect 205140 20480 205360 20520
rect 205140 20410 205150 20480
rect 205350 20410 205360 20480
rect 205140 20360 205360 20410
rect 205640 20590 205860 20640
rect 205640 20520 205650 20590
rect 205850 20520 205860 20590
rect 205640 20480 205860 20520
rect 205640 20410 205650 20480
rect 205850 20410 205860 20480
rect 205640 20360 205860 20410
rect 206140 20590 206360 20640
rect 206140 20520 206150 20590
rect 206350 20520 206360 20590
rect 206140 20480 206360 20520
rect 206140 20410 206150 20480
rect 206350 20410 206360 20480
rect 206140 20360 206360 20410
rect 206640 20590 206860 20640
rect 206640 20520 206650 20590
rect 206850 20520 206860 20590
rect 206640 20480 206860 20520
rect 206640 20410 206650 20480
rect 206850 20410 206860 20480
rect 206640 20360 206860 20410
rect 207140 20590 207360 20640
rect 207140 20520 207150 20590
rect 207350 20520 207360 20590
rect 207140 20480 207360 20520
rect 207140 20410 207150 20480
rect 207350 20410 207360 20480
rect 207140 20360 207360 20410
rect 207640 20590 207860 20640
rect 207640 20520 207650 20590
rect 207850 20520 207860 20590
rect 207640 20480 207860 20520
rect 207640 20410 207650 20480
rect 207850 20410 207860 20480
rect 207640 20360 207860 20410
rect 204000 20350 208000 20360
rect 204000 20150 204020 20350
rect 204090 20150 204410 20350
rect 204480 20150 204520 20350
rect 204590 20150 204910 20350
rect 204980 20150 205020 20350
rect 205090 20150 205410 20350
rect 205480 20150 205520 20350
rect 205590 20150 205910 20350
rect 205980 20150 206020 20350
rect 206090 20150 206410 20350
rect 206480 20150 206520 20350
rect 206590 20150 206910 20350
rect 206980 20150 207020 20350
rect 207090 20150 207410 20350
rect 207480 20150 207520 20350
rect 207590 20150 207910 20350
rect 207980 20150 208000 20350
rect 204000 20140 208000 20150
rect 204140 20090 204360 20140
rect 204140 20020 204150 20090
rect 204350 20020 204360 20090
rect 204140 19980 204360 20020
rect 204140 19910 204150 19980
rect 204350 19910 204360 19980
rect 204140 19860 204360 19910
rect 204640 20090 204860 20140
rect 204640 20020 204650 20090
rect 204850 20020 204860 20090
rect 204640 19980 204860 20020
rect 204640 19910 204650 19980
rect 204850 19910 204860 19980
rect 204640 19860 204860 19910
rect 205140 20090 205360 20140
rect 205140 20020 205150 20090
rect 205350 20020 205360 20090
rect 205140 19980 205360 20020
rect 205140 19910 205150 19980
rect 205350 19910 205360 19980
rect 205140 19860 205360 19910
rect 205640 20090 205860 20140
rect 205640 20020 205650 20090
rect 205850 20020 205860 20090
rect 205640 19980 205860 20020
rect 205640 19910 205650 19980
rect 205850 19910 205860 19980
rect 205640 19860 205860 19910
rect 206140 20090 206360 20140
rect 206140 20020 206150 20090
rect 206350 20020 206360 20090
rect 206140 19980 206360 20020
rect 206140 19910 206150 19980
rect 206350 19910 206360 19980
rect 206140 19860 206360 19910
rect 206640 20090 206860 20140
rect 206640 20020 206650 20090
rect 206850 20020 206860 20090
rect 206640 19980 206860 20020
rect 206640 19910 206650 19980
rect 206850 19910 206860 19980
rect 206640 19860 206860 19910
rect 207140 20090 207360 20140
rect 207140 20020 207150 20090
rect 207350 20020 207360 20090
rect 207140 19980 207360 20020
rect 207140 19910 207150 19980
rect 207350 19910 207360 19980
rect 207140 19860 207360 19910
rect 207640 20090 207860 20140
rect 207640 20020 207650 20090
rect 207850 20020 207860 20090
rect 207640 19980 207860 20020
rect 207640 19910 207650 19980
rect 207850 19910 207860 19980
rect 207640 19860 207860 19910
rect 204000 19850 208000 19860
rect 204000 19650 204020 19850
rect 204090 19650 204410 19850
rect 204480 19650 204520 19850
rect 204590 19650 204910 19850
rect 204980 19650 205020 19850
rect 205090 19650 205410 19850
rect 205480 19650 205520 19850
rect 205590 19650 205910 19850
rect 205980 19650 206020 19850
rect 206090 19650 206410 19850
rect 206480 19650 206520 19850
rect 206590 19650 206910 19850
rect 206980 19650 207020 19850
rect 207090 19650 207410 19850
rect 207480 19650 207520 19850
rect 207590 19650 207910 19850
rect 207980 19650 208000 19850
rect 204000 19640 208000 19650
rect 204140 19590 204360 19640
rect 204140 19520 204150 19590
rect 204350 19520 204360 19590
rect 204140 19480 204360 19520
rect 204140 19410 204150 19480
rect 204350 19410 204360 19480
rect 204140 19360 204360 19410
rect 204640 19590 204860 19640
rect 204640 19520 204650 19590
rect 204850 19520 204860 19590
rect 204640 19480 204860 19520
rect 204640 19410 204650 19480
rect 204850 19410 204860 19480
rect 204640 19360 204860 19410
rect 205140 19590 205360 19640
rect 205140 19520 205150 19590
rect 205350 19520 205360 19590
rect 205140 19480 205360 19520
rect 205140 19410 205150 19480
rect 205350 19410 205360 19480
rect 205140 19360 205360 19410
rect 205640 19590 205860 19640
rect 205640 19520 205650 19590
rect 205850 19520 205860 19590
rect 205640 19480 205860 19520
rect 205640 19410 205650 19480
rect 205850 19410 205860 19480
rect 205640 19360 205860 19410
rect 206140 19590 206360 19640
rect 206140 19520 206150 19590
rect 206350 19520 206360 19590
rect 206140 19480 206360 19520
rect 206140 19410 206150 19480
rect 206350 19410 206360 19480
rect 206140 19360 206360 19410
rect 206640 19590 206860 19640
rect 206640 19520 206650 19590
rect 206850 19520 206860 19590
rect 206640 19480 206860 19520
rect 206640 19410 206650 19480
rect 206850 19410 206860 19480
rect 206640 19360 206860 19410
rect 207140 19590 207360 19640
rect 207140 19520 207150 19590
rect 207350 19520 207360 19590
rect 207140 19480 207360 19520
rect 207140 19410 207150 19480
rect 207350 19410 207360 19480
rect 207140 19360 207360 19410
rect 207640 19590 207860 19640
rect 207640 19520 207650 19590
rect 207850 19520 207860 19590
rect 207640 19480 207860 19520
rect 207640 19410 207650 19480
rect 207850 19410 207860 19480
rect 207640 19360 207860 19410
rect 204000 19350 208000 19360
rect 204000 19150 204020 19350
rect 204090 19150 204410 19350
rect 204480 19150 204520 19350
rect 204590 19150 204910 19350
rect 204980 19150 205020 19350
rect 205090 19150 205410 19350
rect 205480 19150 205520 19350
rect 205590 19150 205910 19350
rect 205980 19150 206020 19350
rect 206090 19150 206410 19350
rect 206480 19150 206520 19350
rect 206590 19150 206910 19350
rect 206980 19150 207020 19350
rect 207090 19150 207410 19350
rect 207480 19150 207520 19350
rect 207590 19150 207910 19350
rect 207980 19150 208000 19350
rect 204000 19140 208000 19150
rect 204140 19090 204360 19140
rect 204140 19020 204150 19090
rect 204350 19020 204360 19090
rect 204140 18980 204360 19020
rect 204140 18910 204150 18980
rect 204350 18910 204360 18980
rect 204140 18860 204360 18910
rect 204640 19090 204860 19140
rect 204640 19020 204650 19090
rect 204850 19020 204860 19090
rect 204640 18980 204860 19020
rect 204640 18910 204650 18980
rect 204850 18910 204860 18980
rect 204640 18860 204860 18910
rect 205140 19090 205360 19140
rect 205140 19020 205150 19090
rect 205350 19020 205360 19090
rect 205140 18980 205360 19020
rect 205140 18910 205150 18980
rect 205350 18910 205360 18980
rect 205140 18860 205360 18910
rect 205640 19090 205860 19140
rect 205640 19020 205650 19090
rect 205850 19020 205860 19090
rect 205640 18980 205860 19020
rect 205640 18910 205650 18980
rect 205850 18910 205860 18980
rect 205640 18860 205860 18910
rect 206140 19090 206360 19140
rect 206140 19020 206150 19090
rect 206350 19020 206360 19090
rect 206140 18980 206360 19020
rect 206140 18910 206150 18980
rect 206350 18910 206360 18980
rect 206140 18860 206360 18910
rect 206640 19090 206860 19140
rect 206640 19020 206650 19090
rect 206850 19020 206860 19090
rect 206640 18980 206860 19020
rect 206640 18910 206650 18980
rect 206850 18910 206860 18980
rect 206640 18860 206860 18910
rect 207140 19090 207360 19140
rect 207140 19020 207150 19090
rect 207350 19020 207360 19090
rect 207140 18980 207360 19020
rect 207140 18910 207150 18980
rect 207350 18910 207360 18980
rect 207140 18860 207360 18910
rect 207640 19090 207860 19140
rect 207640 19020 207650 19090
rect 207850 19020 207860 19090
rect 207640 18980 207860 19020
rect 207640 18910 207650 18980
rect 207850 18910 207860 18980
rect 207640 18860 207860 18910
rect 204000 18850 208000 18860
rect 204000 18650 204020 18850
rect 204090 18650 204410 18850
rect 204480 18650 204520 18850
rect 204590 18650 204910 18850
rect 204980 18650 205020 18850
rect 205090 18650 205410 18850
rect 205480 18650 205520 18850
rect 205590 18650 205910 18850
rect 205980 18650 206020 18850
rect 206090 18650 206410 18850
rect 206480 18650 206520 18850
rect 206590 18650 206910 18850
rect 206980 18650 207020 18850
rect 207090 18650 207410 18850
rect 207480 18650 207520 18850
rect 207590 18650 207910 18850
rect 207980 18650 208000 18850
rect 204000 18640 208000 18650
rect 204140 18590 204360 18640
rect 204140 18520 204150 18590
rect 204350 18520 204360 18590
rect 204140 18480 204360 18520
rect 204140 18410 204150 18480
rect 204350 18410 204360 18480
rect 204140 18360 204360 18410
rect 204640 18590 204860 18640
rect 204640 18520 204650 18590
rect 204850 18520 204860 18590
rect 204640 18480 204860 18520
rect 204640 18410 204650 18480
rect 204850 18410 204860 18480
rect 204640 18360 204860 18410
rect 205140 18590 205360 18640
rect 205140 18520 205150 18590
rect 205350 18520 205360 18590
rect 205140 18480 205360 18520
rect 205140 18410 205150 18480
rect 205350 18410 205360 18480
rect 205140 18360 205360 18410
rect 205640 18590 205860 18640
rect 205640 18520 205650 18590
rect 205850 18520 205860 18590
rect 205640 18480 205860 18520
rect 205640 18410 205650 18480
rect 205850 18410 205860 18480
rect 205640 18360 205860 18410
rect 206140 18590 206360 18640
rect 206140 18520 206150 18590
rect 206350 18520 206360 18590
rect 206140 18480 206360 18520
rect 206140 18410 206150 18480
rect 206350 18410 206360 18480
rect 206140 18360 206360 18410
rect 206640 18590 206860 18640
rect 206640 18520 206650 18590
rect 206850 18520 206860 18590
rect 206640 18480 206860 18520
rect 206640 18410 206650 18480
rect 206850 18410 206860 18480
rect 206640 18360 206860 18410
rect 207140 18590 207360 18640
rect 207140 18520 207150 18590
rect 207350 18520 207360 18590
rect 207140 18480 207360 18520
rect 207140 18410 207150 18480
rect 207350 18410 207360 18480
rect 207140 18360 207360 18410
rect 207640 18590 207860 18640
rect 207640 18520 207650 18590
rect 207850 18520 207860 18590
rect 207640 18480 207860 18520
rect 207640 18410 207650 18480
rect 207850 18410 207860 18480
rect 207640 18360 207860 18410
rect 204000 18350 208000 18360
rect 204000 18150 204020 18350
rect 204090 18150 204410 18350
rect 204480 18150 204520 18350
rect 204590 18150 204910 18350
rect 204980 18150 205020 18350
rect 205090 18150 205410 18350
rect 205480 18150 205520 18350
rect 205590 18150 205910 18350
rect 205980 18150 206020 18350
rect 206090 18150 206410 18350
rect 206480 18150 206520 18350
rect 206590 18150 206910 18350
rect 206980 18150 207020 18350
rect 207090 18150 207410 18350
rect 207480 18150 207520 18350
rect 207590 18150 207910 18350
rect 207980 18150 208000 18350
rect 204000 18140 208000 18150
rect 204140 18090 204360 18140
rect 204140 18020 204150 18090
rect 204350 18020 204360 18090
rect 204140 17980 204360 18020
rect 204140 17910 204150 17980
rect 204350 17910 204360 17980
rect 204140 17860 204360 17910
rect 204640 18090 204860 18140
rect 204640 18020 204650 18090
rect 204850 18020 204860 18090
rect 204640 17980 204860 18020
rect 204640 17910 204650 17980
rect 204850 17910 204860 17980
rect 204640 17860 204860 17910
rect 205140 18090 205360 18140
rect 205140 18020 205150 18090
rect 205350 18020 205360 18090
rect 205140 17980 205360 18020
rect 205140 17910 205150 17980
rect 205350 17910 205360 17980
rect 205140 17860 205360 17910
rect 205640 18090 205860 18140
rect 205640 18020 205650 18090
rect 205850 18020 205860 18090
rect 205640 17980 205860 18020
rect 205640 17910 205650 17980
rect 205850 17910 205860 17980
rect 205640 17860 205860 17910
rect 206140 18090 206360 18140
rect 206140 18020 206150 18090
rect 206350 18020 206360 18090
rect 206140 17980 206360 18020
rect 206140 17910 206150 17980
rect 206350 17910 206360 17980
rect 206140 17860 206360 17910
rect 206640 18090 206860 18140
rect 206640 18020 206650 18090
rect 206850 18020 206860 18090
rect 206640 17980 206860 18020
rect 206640 17910 206650 17980
rect 206850 17910 206860 17980
rect 206640 17860 206860 17910
rect 207140 18090 207360 18140
rect 207140 18020 207150 18090
rect 207350 18020 207360 18090
rect 207140 17980 207360 18020
rect 207140 17910 207150 17980
rect 207350 17910 207360 17980
rect 207140 17860 207360 17910
rect 207640 18090 207860 18140
rect 207640 18020 207650 18090
rect 207850 18020 207860 18090
rect 207640 17980 207860 18020
rect 207640 17910 207650 17980
rect 207850 17910 207860 17980
rect 207640 17860 207860 17910
rect 204000 17850 208000 17860
rect 204000 17650 204020 17850
rect 204090 17650 204410 17850
rect 204480 17650 204520 17850
rect 204590 17650 204910 17850
rect 204980 17650 205020 17850
rect 205090 17650 205410 17850
rect 205480 17650 205520 17850
rect 205590 17650 205910 17850
rect 205980 17650 206020 17850
rect 206090 17650 206410 17850
rect 206480 17650 206520 17850
rect 206590 17650 206910 17850
rect 206980 17650 207020 17850
rect 207090 17650 207410 17850
rect 207480 17650 207520 17850
rect 207590 17650 207910 17850
rect 207980 17650 208000 17850
rect 204000 17640 208000 17650
rect 204140 17590 204360 17640
rect 204140 17520 204150 17590
rect 204350 17520 204360 17590
rect 204140 17480 204360 17520
rect 204140 17410 204150 17480
rect 204350 17410 204360 17480
rect 204140 17360 204360 17410
rect 204640 17590 204860 17640
rect 204640 17520 204650 17590
rect 204850 17520 204860 17590
rect 204640 17480 204860 17520
rect 204640 17410 204650 17480
rect 204850 17410 204860 17480
rect 204640 17360 204860 17410
rect 205140 17590 205360 17640
rect 205140 17520 205150 17590
rect 205350 17520 205360 17590
rect 205140 17480 205360 17520
rect 205140 17410 205150 17480
rect 205350 17410 205360 17480
rect 205140 17360 205360 17410
rect 205640 17590 205860 17640
rect 205640 17520 205650 17590
rect 205850 17520 205860 17590
rect 205640 17480 205860 17520
rect 205640 17410 205650 17480
rect 205850 17410 205860 17480
rect 205640 17360 205860 17410
rect 206140 17590 206360 17640
rect 206140 17520 206150 17590
rect 206350 17520 206360 17590
rect 206140 17480 206360 17520
rect 206140 17410 206150 17480
rect 206350 17410 206360 17480
rect 206140 17360 206360 17410
rect 206640 17590 206860 17640
rect 206640 17520 206650 17590
rect 206850 17520 206860 17590
rect 206640 17480 206860 17520
rect 206640 17410 206650 17480
rect 206850 17410 206860 17480
rect 206640 17360 206860 17410
rect 207140 17590 207360 17640
rect 207140 17520 207150 17590
rect 207350 17520 207360 17590
rect 207140 17480 207360 17520
rect 207140 17410 207150 17480
rect 207350 17410 207360 17480
rect 207140 17360 207360 17410
rect 207640 17590 207860 17640
rect 207640 17520 207650 17590
rect 207850 17520 207860 17590
rect 207640 17480 207860 17520
rect 207640 17410 207650 17480
rect 207850 17410 207860 17480
rect 207640 17360 207860 17410
rect 204000 17350 208000 17360
rect 204000 17150 204020 17350
rect 204090 17150 204410 17350
rect 204480 17150 204520 17350
rect 204590 17150 204910 17350
rect 204980 17150 205020 17350
rect 205090 17150 205410 17350
rect 205480 17150 205520 17350
rect 205590 17150 205910 17350
rect 205980 17150 206020 17350
rect 206090 17150 206410 17350
rect 206480 17150 206520 17350
rect 206590 17150 206910 17350
rect 206980 17150 207020 17350
rect 207090 17150 207410 17350
rect 207480 17150 207520 17350
rect 207590 17150 207910 17350
rect 207980 17150 208000 17350
rect 204000 17140 208000 17150
rect 204140 17090 204360 17140
rect 204140 17020 204150 17090
rect 204350 17020 204360 17090
rect 204140 16980 204360 17020
rect 204140 16910 204150 16980
rect 204350 16910 204360 16980
rect 204140 16860 204360 16910
rect 204640 17090 204860 17140
rect 204640 17020 204650 17090
rect 204850 17020 204860 17090
rect 204640 16980 204860 17020
rect 204640 16910 204650 16980
rect 204850 16910 204860 16980
rect 204640 16860 204860 16910
rect 205140 17090 205360 17140
rect 205140 17020 205150 17090
rect 205350 17020 205360 17090
rect 205140 16980 205360 17020
rect 205140 16910 205150 16980
rect 205350 16910 205360 16980
rect 205140 16860 205360 16910
rect 205640 17090 205860 17140
rect 205640 17020 205650 17090
rect 205850 17020 205860 17090
rect 205640 16980 205860 17020
rect 205640 16910 205650 16980
rect 205850 16910 205860 16980
rect 205640 16860 205860 16910
rect 206140 17090 206360 17140
rect 206140 17020 206150 17090
rect 206350 17020 206360 17090
rect 206140 16980 206360 17020
rect 206140 16910 206150 16980
rect 206350 16910 206360 16980
rect 206140 16860 206360 16910
rect 206640 17090 206860 17140
rect 206640 17020 206650 17090
rect 206850 17020 206860 17090
rect 206640 16980 206860 17020
rect 206640 16910 206650 16980
rect 206850 16910 206860 16980
rect 206640 16860 206860 16910
rect 207140 17090 207360 17140
rect 207140 17020 207150 17090
rect 207350 17020 207360 17090
rect 207140 16980 207360 17020
rect 207140 16910 207150 16980
rect 207350 16910 207360 16980
rect 207140 16860 207360 16910
rect 207640 17090 207860 17140
rect 207640 17020 207650 17090
rect 207850 17020 207860 17090
rect 207640 16980 207860 17020
rect 207640 16910 207650 16980
rect 207850 16910 207860 16980
rect 207640 16860 207860 16910
rect 204000 16850 208000 16860
rect 204000 16650 204020 16850
rect 204090 16650 204410 16850
rect 204480 16650 204520 16850
rect 204590 16650 204910 16850
rect 204980 16650 205020 16850
rect 205090 16650 205410 16850
rect 205480 16650 205520 16850
rect 205590 16650 205910 16850
rect 205980 16650 206020 16850
rect 206090 16650 206410 16850
rect 206480 16650 206520 16850
rect 206590 16650 206910 16850
rect 206980 16650 207020 16850
rect 207090 16650 207410 16850
rect 207480 16650 207520 16850
rect 207590 16650 207910 16850
rect 207980 16650 208000 16850
rect 204000 16640 208000 16650
rect 204140 16590 204360 16640
rect 204140 16520 204150 16590
rect 204350 16520 204360 16590
rect 204140 16480 204360 16520
rect 204140 16410 204150 16480
rect 204350 16410 204360 16480
rect 204140 16360 204360 16410
rect 204640 16590 204860 16640
rect 204640 16520 204650 16590
rect 204850 16520 204860 16590
rect 204640 16480 204860 16520
rect 204640 16410 204650 16480
rect 204850 16410 204860 16480
rect 204640 16360 204860 16410
rect 205140 16590 205360 16640
rect 205140 16520 205150 16590
rect 205350 16520 205360 16590
rect 205140 16480 205360 16520
rect 205140 16410 205150 16480
rect 205350 16410 205360 16480
rect 205140 16360 205360 16410
rect 205640 16590 205860 16640
rect 205640 16520 205650 16590
rect 205850 16520 205860 16590
rect 205640 16480 205860 16520
rect 205640 16410 205650 16480
rect 205850 16410 205860 16480
rect 205640 16360 205860 16410
rect 206140 16590 206360 16640
rect 206140 16520 206150 16590
rect 206350 16520 206360 16590
rect 206140 16480 206360 16520
rect 206140 16410 206150 16480
rect 206350 16410 206360 16480
rect 206140 16360 206360 16410
rect 206640 16590 206860 16640
rect 206640 16520 206650 16590
rect 206850 16520 206860 16590
rect 206640 16480 206860 16520
rect 206640 16410 206650 16480
rect 206850 16410 206860 16480
rect 206640 16360 206860 16410
rect 207140 16590 207360 16640
rect 207140 16520 207150 16590
rect 207350 16520 207360 16590
rect 207140 16480 207360 16520
rect 207140 16410 207150 16480
rect 207350 16410 207360 16480
rect 207140 16360 207360 16410
rect 207640 16590 207860 16640
rect 207640 16520 207650 16590
rect 207850 16520 207860 16590
rect 207640 16480 207860 16520
rect 207640 16410 207650 16480
rect 207850 16410 207860 16480
rect 207640 16360 207860 16410
rect 204000 16350 208000 16360
rect 204000 16150 204020 16350
rect 204090 16150 204410 16350
rect 204480 16150 204520 16350
rect 204590 16150 204910 16350
rect 204980 16150 205020 16350
rect 205090 16150 205410 16350
rect 205480 16150 205520 16350
rect 205590 16150 205910 16350
rect 205980 16150 206020 16350
rect 206090 16150 206410 16350
rect 206480 16150 206520 16350
rect 206590 16150 206910 16350
rect 206980 16150 207020 16350
rect 207090 16150 207410 16350
rect 207480 16150 207520 16350
rect 207590 16150 207910 16350
rect 207980 16150 208000 16350
rect 204000 16140 208000 16150
rect 204140 16090 204360 16140
rect 204140 16020 204150 16090
rect 204350 16020 204360 16090
rect 204140 15980 204360 16020
rect 204140 15910 204150 15980
rect 204350 15910 204360 15980
rect 204140 15860 204360 15910
rect 204640 16090 204860 16140
rect 204640 16020 204650 16090
rect 204850 16020 204860 16090
rect 204640 15980 204860 16020
rect 204640 15910 204650 15980
rect 204850 15910 204860 15980
rect 204640 15860 204860 15910
rect 205140 16090 205360 16140
rect 205140 16020 205150 16090
rect 205350 16020 205360 16090
rect 205140 15980 205360 16020
rect 205140 15910 205150 15980
rect 205350 15910 205360 15980
rect 205140 15860 205360 15910
rect 205640 16090 205860 16140
rect 205640 16020 205650 16090
rect 205850 16020 205860 16090
rect 205640 15980 205860 16020
rect 205640 15910 205650 15980
rect 205850 15910 205860 15980
rect 205640 15860 205860 15910
rect 206140 16090 206360 16140
rect 206140 16020 206150 16090
rect 206350 16020 206360 16090
rect 206140 15980 206360 16020
rect 206140 15910 206150 15980
rect 206350 15910 206360 15980
rect 206140 15860 206360 15910
rect 206640 16090 206860 16140
rect 206640 16020 206650 16090
rect 206850 16020 206860 16090
rect 206640 15980 206860 16020
rect 206640 15910 206650 15980
rect 206850 15910 206860 15980
rect 206640 15860 206860 15910
rect 207140 16090 207360 16140
rect 207140 16020 207150 16090
rect 207350 16020 207360 16090
rect 207140 15980 207360 16020
rect 207140 15910 207150 15980
rect 207350 15910 207360 15980
rect 207140 15860 207360 15910
rect 207640 16090 207860 16140
rect 207640 16020 207650 16090
rect 207850 16020 207860 16090
rect 207640 15980 207860 16020
rect 207640 15910 207650 15980
rect 207850 15910 207860 15980
rect 207640 15860 207860 15910
rect 204000 15850 208000 15860
rect 204000 15650 204020 15850
rect 204090 15650 204410 15850
rect 204480 15650 204520 15850
rect 204590 15650 204910 15850
rect 204980 15650 205020 15850
rect 205090 15650 205410 15850
rect 205480 15650 205520 15850
rect 205590 15650 205910 15850
rect 205980 15650 206020 15850
rect 206090 15650 206410 15850
rect 206480 15650 206520 15850
rect 206590 15650 206910 15850
rect 206980 15650 207020 15850
rect 207090 15650 207410 15850
rect 207480 15650 207520 15850
rect 207590 15650 207910 15850
rect 207980 15650 208000 15850
rect 204000 15640 208000 15650
rect 204140 15590 204360 15640
rect 204140 15520 204150 15590
rect 204350 15520 204360 15590
rect 204140 15480 204360 15520
rect 204140 15410 204150 15480
rect 204350 15410 204360 15480
rect 204140 15360 204360 15410
rect 204640 15590 204860 15640
rect 204640 15520 204650 15590
rect 204850 15520 204860 15590
rect 204640 15480 204860 15520
rect 204640 15410 204650 15480
rect 204850 15410 204860 15480
rect 204640 15360 204860 15410
rect 205140 15590 205360 15640
rect 205140 15520 205150 15590
rect 205350 15520 205360 15590
rect 205140 15480 205360 15520
rect 205140 15410 205150 15480
rect 205350 15410 205360 15480
rect 205140 15360 205360 15410
rect 205640 15590 205860 15640
rect 205640 15520 205650 15590
rect 205850 15520 205860 15590
rect 205640 15480 205860 15520
rect 205640 15410 205650 15480
rect 205850 15410 205860 15480
rect 205640 15360 205860 15410
rect 206140 15590 206360 15640
rect 206140 15520 206150 15590
rect 206350 15520 206360 15590
rect 206140 15480 206360 15520
rect 206140 15410 206150 15480
rect 206350 15410 206360 15480
rect 206140 15360 206360 15410
rect 206640 15590 206860 15640
rect 206640 15520 206650 15590
rect 206850 15520 206860 15590
rect 206640 15480 206860 15520
rect 206640 15410 206650 15480
rect 206850 15410 206860 15480
rect 206640 15360 206860 15410
rect 207140 15590 207360 15640
rect 207140 15520 207150 15590
rect 207350 15520 207360 15590
rect 207140 15480 207360 15520
rect 207140 15410 207150 15480
rect 207350 15410 207360 15480
rect 207140 15360 207360 15410
rect 207640 15590 207860 15640
rect 207640 15520 207650 15590
rect 207850 15520 207860 15590
rect 207640 15480 207860 15520
rect 207640 15410 207650 15480
rect 207850 15410 207860 15480
rect 207640 15360 207860 15410
rect 204000 15350 208000 15360
rect 204000 15150 204020 15350
rect 204090 15150 204410 15350
rect 204480 15150 204520 15350
rect 204590 15150 204910 15350
rect 204980 15150 205020 15350
rect 205090 15150 205410 15350
rect 205480 15150 205520 15350
rect 205590 15150 205910 15350
rect 205980 15150 206020 15350
rect 206090 15150 206410 15350
rect 206480 15150 206520 15350
rect 206590 15150 206910 15350
rect 206980 15150 207020 15350
rect 207090 15150 207410 15350
rect 207480 15150 207520 15350
rect 207590 15150 207910 15350
rect 207980 15150 208000 15350
rect 204000 15140 208000 15150
rect 204140 15090 204360 15140
rect 204140 15020 204150 15090
rect 204350 15020 204360 15090
rect 204140 14980 204360 15020
rect 204140 14910 204150 14980
rect 204350 14910 204360 14980
rect 204140 14860 204360 14910
rect 204640 15090 204860 15140
rect 204640 15020 204650 15090
rect 204850 15020 204860 15090
rect 204640 14980 204860 15020
rect 204640 14910 204650 14980
rect 204850 14910 204860 14980
rect 204640 14860 204860 14910
rect 205140 15090 205360 15140
rect 205140 15020 205150 15090
rect 205350 15020 205360 15090
rect 205140 14980 205360 15020
rect 205140 14910 205150 14980
rect 205350 14910 205360 14980
rect 205140 14860 205360 14910
rect 205640 15090 205860 15140
rect 205640 15020 205650 15090
rect 205850 15020 205860 15090
rect 205640 14980 205860 15020
rect 205640 14910 205650 14980
rect 205850 14910 205860 14980
rect 205640 14860 205860 14910
rect 206140 15090 206360 15140
rect 206140 15020 206150 15090
rect 206350 15020 206360 15090
rect 206140 14980 206360 15020
rect 206140 14910 206150 14980
rect 206350 14910 206360 14980
rect 206140 14860 206360 14910
rect 206640 15090 206860 15140
rect 206640 15020 206650 15090
rect 206850 15020 206860 15090
rect 206640 14980 206860 15020
rect 206640 14910 206650 14980
rect 206850 14910 206860 14980
rect 206640 14860 206860 14910
rect 207140 15090 207360 15140
rect 207140 15020 207150 15090
rect 207350 15020 207360 15090
rect 207140 14980 207360 15020
rect 207140 14910 207150 14980
rect 207350 14910 207360 14980
rect 207140 14860 207360 14910
rect 207640 15090 207860 15140
rect 207640 15020 207650 15090
rect 207850 15020 207860 15090
rect 207640 14980 207860 15020
rect 207640 14910 207650 14980
rect 207850 14910 207860 14980
rect 207640 14860 207860 14910
rect 204000 14850 208000 14860
rect 204000 14650 204020 14850
rect 204090 14650 204410 14850
rect 204480 14650 204520 14850
rect 204590 14650 204910 14850
rect 204980 14650 205020 14850
rect 205090 14650 205410 14850
rect 205480 14650 205520 14850
rect 205590 14650 205910 14850
rect 205980 14650 206020 14850
rect 206090 14650 206410 14850
rect 206480 14650 206520 14850
rect 206590 14650 206910 14850
rect 206980 14650 207020 14850
rect 207090 14650 207410 14850
rect 207480 14650 207520 14850
rect 207590 14650 207910 14850
rect 207980 14650 208000 14850
rect 204000 14640 208000 14650
rect 204140 14590 204360 14640
rect 204140 14520 204150 14590
rect 204350 14520 204360 14590
rect 204140 14480 204360 14520
rect 204140 14410 204150 14480
rect 204350 14410 204360 14480
rect 204140 14360 204360 14410
rect 204640 14590 204860 14640
rect 204640 14520 204650 14590
rect 204850 14520 204860 14590
rect 204640 14480 204860 14520
rect 204640 14410 204650 14480
rect 204850 14410 204860 14480
rect 204640 14360 204860 14410
rect 205140 14590 205360 14640
rect 205140 14520 205150 14590
rect 205350 14520 205360 14590
rect 205140 14480 205360 14520
rect 205140 14410 205150 14480
rect 205350 14410 205360 14480
rect 205140 14360 205360 14410
rect 205640 14590 205860 14640
rect 205640 14520 205650 14590
rect 205850 14520 205860 14590
rect 205640 14480 205860 14520
rect 205640 14410 205650 14480
rect 205850 14410 205860 14480
rect 205640 14360 205860 14410
rect 206140 14590 206360 14640
rect 206140 14520 206150 14590
rect 206350 14520 206360 14590
rect 206140 14480 206360 14520
rect 206140 14410 206150 14480
rect 206350 14410 206360 14480
rect 206140 14360 206360 14410
rect 206640 14590 206860 14640
rect 206640 14520 206650 14590
rect 206850 14520 206860 14590
rect 206640 14480 206860 14520
rect 206640 14410 206650 14480
rect 206850 14410 206860 14480
rect 206640 14360 206860 14410
rect 207140 14590 207360 14640
rect 207140 14520 207150 14590
rect 207350 14520 207360 14590
rect 207140 14480 207360 14520
rect 207140 14410 207150 14480
rect 207350 14410 207360 14480
rect 207140 14360 207360 14410
rect 207640 14590 207860 14640
rect 207640 14520 207650 14590
rect 207850 14520 207860 14590
rect 207640 14480 207860 14520
rect 207640 14410 207650 14480
rect 207850 14410 207860 14480
rect 207640 14360 207860 14410
rect 204000 14350 208000 14360
rect 204000 14150 204020 14350
rect 204090 14150 204410 14350
rect 204480 14150 204520 14350
rect 204590 14150 204910 14350
rect 204980 14150 205020 14350
rect 205090 14150 205410 14350
rect 205480 14150 205520 14350
rect 205590 14150 205910 14350
rect 205980 14150 206020 14350
rect 206090 14150 206410 14350
rect 206480 14150 206520 14350
rect 206590 14150 206910 14350
rect 206980 14150 207020 14350
rect 207090 14150 207410 14350
rect 207480 14150 207520 14350
rect 207590 14150 207910 14350
rect 207980 14150 208000 14350
rect 204000 14140 208000 14150
rect 204140 14090 204360 14140
rect 204140 14020 204150 14090
rect 204350 14020 204360 14090
rect 204140 13980 204360 14020
rect 204140 13910 204150 13980
rect 204350 13910 204360 13980
rect 204140 13860 204360 13910
rect 204640 14090 204860 14140
rect 204640 14020 204650 14090
rect 204850 14020 204860 14090
rect 204640 13980 204860 14020
rect 204640 13910 204650 13980
rect 204850 13910 204860 13980
rect 204640 13860 204860 13910
rect 205140 14090 205360 14140
rect 205140 14020 205150 14090
rect 205350 14020 205360 14090
rect 205140 13980 205360 14020
rect 205140 13910 205150 13980
rect 205350 13910 205360 13980
rect 205140 13860 205360 13910
rect 205640 14090 205860 14140
rect 205640 14020 205650 14090
rect 205850 14020 205860 14090
rect 205640 13980 205860 14020
rect 205640 13910 205650 13980
rect 205850 13910 205860 13980
rect 205640 13860 205860 13910
rect 206140 14090 206360 14140
rect 206140 14020 206150 14090
rect 206350 14020 206360 14090
rect 206140 13980 206360 14020
rect 206140 13910 206150 13980
rect 206350 13910 206360 13980
rect 206140 13860 206360 13910
rect 206640 14090 206860 14140
rect 206640 14020 206650 14090
rect 206850 14020 206860 14090
rect 206640 13980 206860 14020
rect 206640 13910 206650 13980
rect 206850 13910 206860 13980
rect 206640 13860 206860 13910
rect 207140 14090 207360 14140
rect 207140 14020 207150 14090
rect 207350 14020 207360 14090
rect 207140 13980 207360 14020
rect 207140 13910 207150 13980
rect 207350 13910 207360 13980
rect 207140 13860 207360 13910
rect 207640 14090 207860 14140
rect 207640 14020 207650 14090
rect 207850 14020 207860 14090
rect 207640 13980 207860 14020
rect 207640 13910 207650 13980
rect 207850 13910 207860 13980
rect 207640 13860 207860 13910
rect 204000 13850 208000 13860
rect 204000 13650 204020 13850
rect 204090 13650 204410 13850
rect 204480 13650 204520 13850
rect 204590 13650 204910 13850
rect 204980 13650 205020 13850
rect 205090 13650 205410 13850
rect 205480 13650 205520 13850
rect 205590 13650 205910 13850
rect 205980 13650 206020 13850
rect 206090 13650 206410 13850
rect 206480 13650 206520 13850
rect 206590 13650 206910 13850
rect 206980 13650 207020 13850
rect 207090 13650 207410 13850
rect 207480 13650 207520 13850
rect 207590 13650 207910 13850
rect 207980 13650 208000 13850
rect 204000 13640 208000 13650
rect 204140 13590 204360 13640
rect 204140 13520 204150 13590
rect 204350 13520 204360 13590
rect 204140 13480 204360 13520
rect 204140 13410 204150 13480
rect 204350 13410 204360 13480
rect 204140 13360 204360 13410
rect 204640 13590 204860 13640
rect 204640 13520 204650 13590
rect 204850 13520 204860 13590
rect 204640 13480 204860 13520
rect 204640 13410 204650 13480
rect 204850 13410 204860 13480
rect 204640 13360 204860 13410
rect 205140 13590 205360 13640
rect 205140 13520 205150 13590
rect 205350 13520 205360 13590
rect 205140 13480 205360 13520
rect 205140 13410 205150 13480
rect 205350 13410 205360 13480
rect 205140 13360 205360 13410
rect 205640 13590 205860 13640
rect 205640 13520 205650 13590
rect 205850 13520 205860 13590
rect 205640 13480 205860 13520
rect 205640 13410 205650 13480
rect 205850 13410 205860 13480
rect 205640 13360 205860 13410
rect 206140 13590 206360 13640
rect 206140 13520 206150 13590
rect 206350 13520 206360 13590
rect 206140 13480 206360 13520
rect 206140 13410 206150 13480
rect 206350 13410 206360 13480
rect 206140 13360 206360 13410
rect 206640 13590 206860 13640
rect 206640 13520 206650 13590
rect 206850 13520 206860 13590
rect 206640 13480 206860 13520
rect 206640 13410 206650 13480
rect 206850 13410 206860 13480
rect 206640 13360 206860 13410
rect 207140 13590 207360 13640
rect 207140 13520 207150 13590
rect 207350 13520 207360 13590
rect 207140 13480 207360 13520
rect 207140 13410 207150 13480
rect 207350 13410 207360 13480
rect 207140 13360 207360 13410
rect 207640 13590 207860 13640
rect 207640 13520 207650 13590
rect 207850 13520 207860 13590
rect 207640 13480 207860 13520
rect 207640 13410 207650 13480
rect 207850 13410 207860 13480
rect 207640 13360 207860 13410
rect 204000 13350 208000 13360
rect 204000 13150 204020 13350
rect 204090 13150 204410 13350
rect 204480 13150 204520 13350
rect 204590 13150 204910 13350
rect 204980 13150 205020 13350
rect 205090 13150 205410 13350
rect 205480 13150 205520 13350
rect 205590 13150 205910 13350
rect 205980 13150 206020 13350
rect 206090 13150 206410 13350
rect 206480 13150 206520 13350
rect 206590 13150 206910 13350
rect 206980 13150 207020 13350
rect 207090 13150 207410 13350
rect 207480 13150 207520 13350
rect 207590 13150 207910 13350
rect 207980 13150 208000 13350
rect 204000 13140 208000 13150
rect 204140 13090 204360 13140
rect 204140 13020 204150 13090
rect 204350 13020 204360 13090
rect 204140 12980 204360 13020
rect 204140 12910 204150 12980
rect 204350 12910 204360 12980
rect 204140 12860 204360 12910
rect 204640 13090 204860 13140
rect 204640 13020 204650 13090
rect 204850 13020 204860 13090
rect 204640 12980 204860 13020
rect 204640 12910 204650 12980
rect 204850 12910 204860 12980
rect 204640 12860 204860 12910
rect 205140 13090 205360 13140
rect 205140 13020 205150 13090
rect 205350 13020 205360 13090
rect 205140 12980 205360 13020
rect 205140 12910 205150 12980
rect 205350 12910 205360 12980
rect 205140 12860 205360 12910
rect 205640 13090 205860 13140
rect 205640 13020 205650 13090
rect 205850 13020 205860 13090
rect 205640 12980 205860 13020
rect 205640 12910 205650 12980
rect 205850 12910 205860 12980
rect 205640 12860 205860 12910
rect 206140 13090 206360 13140
rect 206140 13020 206150 13090
rect 206350 13020 206360 13090
rect 206140 12980 206360 13020
rect 206140 12910 206150 12980
rect 206350 12910 206360 12980
rect 206140 12860 206360 12910
rect 206640 13090 206860 13140
rect 206640 13020 206650 13090
rect 206850 13020 206860 13090
rect 206640 12980 206860 13020
rect 206640 12910 206650 12980
rect 206850 12910 206860 12980
rect 206640 12860 206860 12910
rect 207140 13090 207360 13140
rect 207140 13020 207150 13090
rect 207350 13020 207360 13090
rect 207140 12980 207360 13020
rect 207140 12910 207150 12980
rect 207350 12910 207360 12980
rect 207140 12860 207360 12910
rect 207640 13090 207860 13140
rect 207640 13020 207650 13090
rect 207850 13020 207860 13090
rect 207640 12980 207860 13020
rect 207640 12910 207650 12980
rect 207850 12910 207860 12980
rect 207640 12860 207860 12910
rect 204000 12850 208000 12860
rect 204000 12650 204020 12850
rect 204090 12650 204410 12850
rect 204480 12650 204520 12850
rect 204590 12650 204910 12850
rect 204980 12650 205020 12850
rect 205090 12650 205410 12850
rect 205480 12650 205520 12850
rect 205590 12650 205910 12850
rect 205980 12650 206020 12850
rect 206090 12650 206410 12850
rect 206480 12650 206520 12850
rect 206590 12650 206910 12850
rect 206980 12650 207020 12850
rect 207090 12650 207410 12850
rect 207480 12650 207520 12850
rect 207590 12650 207910 12850
rect 207980 12650 208000 12850
rect 204000 12640 208000 12650
rect 204140 12590 204360 12640
rect 204140 12520 204150 12590
rect 204350 12520 204360 12590
rect 204140 12480 204360 12520
rect 204140 12410 204150 12480
rect 204350 12410 204360 12480
rect 204140 12360 204360 12410
rect 204640 12590 204860 12640
rect 204640 12520 204650 12590
rect 204850 12520 204860 12590
rect 204640 12480 204860 12520
rect 204640 12410 204650 12480
rect 204850 12410 204860 12480
rect 204640 12360 204860 12410
rect 205140 12590 205360 12640
rect 205140 12520 205150 12590
rect 205350 12520 205360 12590
rect 205140 12480 205360 12520
rect 205140 12410 205150 12480
rect 205350 12410 205360 12480
rect 205140 12360 205360 12410
rect 205640 12590 205860 12640
rect 205640 12520 205650 12590
rect 205850 12520 205860 12590
rect 205640 12480 205860 12520
rect 205640 12410 205650 12480
rect 205850 12410 205860 12480
rect 205640 12360 205860 12410
rect 206140 12590 206360 12640
rect 206140 12520 206150 12590
rect 206350 12520 206360 12590
rect 206140 12480 206360 12520
rect 206140 12410 206150 12480
rect 206350 12410 206360 12480
rect 206140 12360 206360 12410
rect 206640 12590 206860 12640
rect 206640 12520 206650 12590
rect 206850 12520 206860 12590
rect 206640 12480 206860 12520
rect 206640 12410 206650 12480
rect 206850 12410 206860 12480
rect 206640 12360 206860 12410
rect 207140 12590 207360 12640
rect 207140 12520 207150 12590
rect 207350 12520 207360 12590
rect 207140 12480 207360 12520
rect 207140 12410 207150 12480
rect 207350 12410 207360 12480
rect 207140 12360 207360 12410
rect 207640 12590 207860 12640
rect 207640 12520 207650 12590
rect 207850 12520 207860 12590
rect 207640 12480 207860 12520
rect 207640 12410 207650 12480
rect 207850 12410 207860 12480
rect 207640 12360 207860 12410
rect 204000 12350 208000 12360
rect 204000 12150 204020 12350
rect 204090 12150 204410 12350
rect 204480 12150 204520 12350
rect 204590 12150 204910 12350
rect 204980 12150 205020 12350
rect 205090 12150 205410 12350
rect 205480 12150 205520 12350
rect 205590 12150 205910 12350
rect 205980 12150 206020 12350
rect 206090 12150 206410 12350
rect 206480 12150 206520 12350
rect 206590 12150 206910 12350
rect 206980 12150 207020 12350
rect 207090 12150 207410 12350
rect 207480 12150 207520 12350
rect 207590 12150 207910 12350
rect 207980 12150 208000 12350
rect 204000 12140 208000 12150
rect 204140 12090 204360 12140
rect 204140 12020 204150 12090
rect 204350 12020 204360 12090
rect 204140 11980 204360 12020
rect 204140 11910 204150 11980
rect 204350 11910 204360 11980
rect 204140 11860 204360 11910
rect 204640 12090 204860 12140
rect 204640 12020 204650 12090
rect 204850 12020 204860 12090
rect 204640 11980 204860 12020
rect 204640 11910 204650 11980
rect 204850 11910 204860 11980
rect 204640 11860 204860 11910
rect 205140 12090 205360 12140
rect 205140 12020 205150 12090
rect 205350 12020 205360 12090
rect 205140 11980 205360 12020
rect 205140 11910 205150 11980
rect 205350 11910 205360 11980
rect 205140 11860 205360 11910
rect 205640 12090 205860 12140
rect 205640 12020 205650 12090
rect 205850 12020 205860 12090
rect 205640 11980 205860 12020
rect 205640 11910 205650 11980
rect 205850 11910 205860 11980
rect 205640 11860 205860 11910
rect 206140 12090 206360 12140
rect 206140 12020 206150 12090
rect 206350 12020 206360 12090
rect 206140 11980 206360 12020
rect 206140 11910 206150 11980
rect 206350 11910 206360 11980
rect 206140 11860 206360 11910
rect 206640 12090 206860 12140
rect 206640 12020 206650 12090
rect 206850 12020 206860 12090
rect 206640 11980 206860 12020
rect 206640 11910 206650 11980
rect 206850 11910 206860 11980
rect 206640 11860 206860 11910
rect 207140 12090 207360 12140
rect 207140 12020 207150 12090
rect 207350 12020 207360 12090
rect 207140 11980 207360 12020
rect 207140 11910 207150 11980
rect 207350 11910 207360 11980
rect 207140 11860 207360 11910
rect 207640 12090 207860 12140
rect 207640 12020 207650 12090
rect 207850 12020 207860 12090
rect 207640 11980 207860 12020
rect 207640 11910 207650 11980
rect 207850 11910 207860 11980
rect 207640 11860 207860 11910
rect 204000 11850 208000 11860
rect 204000 11650 204020 11850
rect 204090 11650 204410 11850
rect 204480 11650 204520 11850
rect 204590 11650 204910 11850
rect 204980 11650 205020 11850
rect 205090 11650 205410 11850
rect 205480 11650 205520 11850
rect 205590 11650 205910 11850
rect 205980 11650 206020 11850
rect 206090 11650 206410 11850
rect 206480 11650 206520 11850
rect 206590 11650 206910 11850
rect 206980 11650 207020 11850
rect 207090 11650 207410 11850
rect 207480 11650 207520 11850
rect 207590 11650 207910 11850
rect 207980 11650 208000 11850
rect 204000 11640 208000 11650
rect 204140 11590 204360 11640
rect 204140 11520 204150 11590
rect 204350 11520 204360 11590
rect 204140 11480 204360 11520
rect 204140 11410 204150 11480
rect 204350 11410 204360 11480
rect 204140 11360 204360 11410
rect 204640 11590 204860 11640
rect 204640 11520 204650 11590
rect 204850 11520 204860 11590
rect 204640 11480 204860 11520
rect 204640 11410 204650 11480
rect 204850 11410 204860 11480
rect 204640 11360 204860 11410
rect 205140 11590 205360 11640
rect 205140 11520 205150 11590
rect 205350 11520 205360 11590
rect 205140 11480 205360 11520
rect 205140 11410 205150 11480
rect 205350 11410 205360 11480
rect 205140 11360 205360 11410
rect 205640 11590 205860 11640
rect 205640 11520 205650 11590
rect 205850 11520 205860 11590
rect 205640 11480 205860 11520
rect 205640 11410 205650 11480
rect 205850 11410 205860 11480
rect 205640 11360 205860 11410
rect 206140 11590 206360 11640
rect 206140 11520 206150 11590
rect 206350 11520 206360 11590
rect 206140 11480 206360 11520
rect 206140 11410 206150 11480
rect 206350 11410 206360 11480
rect 206140 11360 206360 11410
rect 206640 11590 206860 11640
rect 206640 11520 206650 11590
rect 206850 11520 206860 11590
rect 206640 11480 206860 11520
rect 206640 11410 206650 11480
rect 206850 11410 206860 11480
rect 206640 11360 206860 11410
rect 207140 11590 207360 11640
rect 207140 11520 207150 11590
rect 207350 11520 207360 11590
rect 207140 11480 207360 11520
rect 207140 11410 207150 11480
rect 207350 11410 207360 11480
rect 207140 11360 207360 11410
rect 207640 11590 207860 11640
rect 207640 11520 207650 11590
rect 207850 11520 207860 11590
rect 207640 11480 207860 11520
rect 207640 11410 207650 11480
rect 207850 11410 207860 11480
rect 207640 11360 207860 11410
rect 204000 11350 208000 11360
rect 204000 11150 204020 11350
rect 204090 11150 204410 11350
rect 204480 11150 204520 11350
rect 204590 11150 204910 11350
rect 204980 11150 205020 11350
rect 205090 11150 205410 11350
rect 205480 11150 205520 11350
rect 205590 11150 205910 11350
rect 205980 11150 206020 11350
rect 206090 11150 206410 11350
rect 206480 11150 206520 11350
rect 206590 11150 206910 11350
rect 206980 11150 207020 11350
rect 207090 11150 207410 11350
rect 207480 11150 207520 11350
rect 207590 11150 207910 11350
rect 207980 11150 208000 11350
rect 204000 11140 208000 11150
rect 204140 11090 204360 11140
rect 204140 11020 204150 11090
rect 204350 11020 204360 11090
rect 204140 10980 204360 11020
rect 204140 10910 204150 10980
rect 204350 10910 204360 10980
rect 204140 10860 204360 10910
rect 204640 11090 204860 11140
rect 204640 11020 204650 11090
rect 204850 11020 204860 11090
rect 204640 10980 204860 11020
rect 204640 10910 204650 10980
rect 204850 10910 204860 10980
rect 204640 10860 204860 10910
rect 205140 11090 205360 11140
rect 205140 11020 205150 11090
rect 205350 11020 205360 11090
rect 205140 10980 205360 11020
rect 205140 10910 205150 10980
rect 205350 10910 205360 10980
rect 205140 10860 205360 10910
rect 205640 11090 205860 11140
rect 205640 11020 205650 11090
rect 205850 11020 205860 11090
rect 205640 10980 205860 11020
rect 205640 10910 205650 10980
rect 205850 10910 205860 10980
rect 205640 10860 205860 10910
rect 206140 11090 206360 11140
rect 206140 11020 206150 11090
rect 206350 11020 206360 11090
rect 206140 10980 206360 11020
rect 206140 10910 206150 10980
rect 206350 10910 206360 10980
rect 206140 10860 206360 10910
rect 206640 11090 206860 11140
rect 206640 11020 206650 11090
rect 206850 11020 206860 11090
rect 206640 10980 206860 11020
rect 206640 10910 206650 10980
rect 206850 10910 206860 10980
rect 206640 10860 206860 10910
rect 207140 11090 207360 11140
rect 207140 11020 207150 11090
rect 207350 11020 207360 11090
rect 207140 10980 207360 11020
rect 207140 10910 207150 10980
rect 207350 10910 207360 10980
rect 207140 10860 207360 10910
rect 207640 11090 207860 11140
rect 207640 11020 207650 11090
rect 207850 11020 207860 11090
rect 207640 10980 207860 11020
rect 207640 10910 207650 10980
rect 207850 10910 207860 10980
rect 207640 10860 207860 10910
rect 204000 10850 208000 10860
rect 204000 10650 204020 10850
rect 204090 10650 204410 10850
rect 204480 10650 204520 10850
rect 204590 10650 204910 10850
rect 204980 10650 205020 10850
rect 205090 10650 205410 10850
rect 205480 10650 205520 10850
rect 205590 10650 205910 10850
rect 205980 10650 206020 10850
rect 206090 10650 206410 10850
rect 206480 10650 206520 10850
rect 206590 10650 206910 10850
rect 206980 10650 207020 10850
rect 207090 10650 207410 10850
rect 207480 10650 207520 10850
rect 207590 10650 207910 10850
rect 207980 10650 208000 10850
rect 204000 10640 208000 10650
rect 204140 10590 204360 10640
rect 204140 10520 204150 10590
rect 204350 10520 204360 10590
rect 204140 10480 204360 10520
rect 204140 10410 204150 10480
rect 204350 10410 204360 10480
rect 204140 10360 204360 10410
rect 204640 10590 204860 10640
rect 204640 10520 204650 10590
rect 204850 10520 204860 10590
rect 204640 10480 204860 10520
rect 204640 10410 204650 10480
rect 204850 10410 204860 10480
rect 204640 10360 204860 10410
rect 205140 10590 205360 10640
rect 205140 10520 205150 10590
rect 205350 10520 205360 10590
rect 205140 10480 205360 10520
rect 205140 10410 205150 10480
rect 205350 10410 205360 10480
rect 205140 10360 205360 10410
rect 205640 10590 205860 10640
rect 205640 10520 205650 10590
rect 205850 10520 205860 10590
rect 205640 10480 205860 10520
rect 205640 10410 205650 10480
rect 205850 10410 205860 10480
rect 205640 10360 205860 10410
rect 206140 10590 206360 10640
rect 206140 10520 206150 10590
rect 206350 10520 206360 10590
rect 206140 10480 206360 10520
rect 206140 10410 206150 10480
rect 206350 10410 206360 10480
rect 206140 10360 206360 10410
rect 206640 10590 206860 10640
rect 206640 10520 206650 10590
rect 206850 10520 206860 10590
rect 206640 10480 206860 10520
rect 206640 10410 206650 10480
rect 206850 10410 206860 10480
rect 206640 10360 206860 10410
rect 207140 10590 207360 10640
rect 207140 10520 207150 10590
rect 207350 10520 207360 10590
rect 207140 10480 207360 10520
rect 207140 10410 207150 10480
rect 207350 10410 207360 10480
rect 207140 10360 207360 10410
rect 207640 10590 207860 10640
rect 207640 10520 207650 10590
rect 207850 10520 207860 10590
rect 207640 10480 207860 10520
rect 207640 10410 207650 10480
rect 207850 10410 207860 10480
rect 207640 10360 207860 10410
rect 204000 10350 208000 10360
rect 204000 10150 204020 10350
rect 204090 10150 204410 10350
rect 204480 10150 204520 10350
rect 204590 10150 204910 10350
rect 204980 10150 205020 10350
rect 205090 10150 205410 10350
rect 205480 10150 205520 10350
rect 205590 10150 205910 10350
rect 205980 10150 206020 10350
rect 206090 10150 206410 10350
rect 206480 10150 206520 10350
rect 206590 10150 206910 10350
rect 206980 10150 207020 10350
rect 207090 10150 207410 10350
rect 207480 10150 207520 10350
rect 207590 10150 207910 10350
rect 207980 10150 208000 10350
rect 204000 10140 208000 10150
rect 204140 10090 204360 10140
rect 204140 10020 204150 10090
rect 204350 10020 204360 10090
rect 204140 9980 204360 10020
rect 204140 9910 204150 9980
rect 204350 9910 204360 9980
rect 204140 9860 204360 9910
rect 204640 10090 204860 10140
rect 204640 10020 204650 10090
rect 204850 10020 204860 10090
rect 204640 9980 204860 10020
rect 204640 9910 204650 9980
rect 204850 9910 204860 9980
rect 204640 9860 204860 9910
rect 205140 10090 205360 10140
rect 205140 10020 205150 10090
rect 205350 10020 205360 10090
rect 205140 9980 205360 10020
rect 205140 9910 205150 9980
rect 205350 9910 205360 9980
rect 205140 9860 205360 9910
rect 205640 10090 205860 10140
rect 205640 10020 205650 10090
rect 205850 10020 205860 10090
rect 205640 9980 205860 10020
rect 205640 9910 205650 9980
rect 205850 9910 205860 9980
rect 205640 9860 205860 9910
rect 206140 10090 206360 10140
rect 206140 10020 206150 10090
rect 206350 10020 206360 10090
rect 206140 9980 206360 10020
rect 206140 9910 206150 9980
rect 206350 9910 206360 9980
rect 206140 9860 206360 9910
rect 206640 10090 206860 10140
rect 206640 10020 206650 10090
rect 206850 10020 206860 10090
rect 206640 9980 206860 10020
rect 206640 9910 206650 9980
rect 206850 9910 206860 9980
rect 206640 9860 206860 9910
rect 207140 10090 207360 10140
rect 207140 10020 207150 10090
rect 207350 10020 207360 10090
rect 207140 9980 207360 10020
rect 207140 9910 207150 9980
rect 207350 9910 207360 9980
rect 207140 9860 207360 9910
rect 207640 10090 207860 10140
rect 207640 10020 207650 10090
rect 207850 10020 207860 10090
rect 207640 9980 207860 10020
rect 207640 9910 207650 9980
rect 207850 9910 207860 9980
rect 207640 9860 207860 9910
rect 204000 9850 208000 9860
rect 204000 9650 204020 9850
rect 204090 9650 204410 9850
rect 204480 9650 204520 9850
rect 204590 9650 204910 9850
rect 204980 9650 205020 9850
rect 205090 9650 205410 9850
rect 205480 9650 205520 9850
rect 205590 9650 205910 9850
rect 205980 9650 206020 9850
rect 206090 9650 206410 9850
rect 206480 9650 206520 9850
rect 206590 9650 206910 9850
rect 206980 9650 207020 9850
rect 207090 9650 207410 9850
rect 207480 9650 207520 9850
rect 207590 9650 207910 9850
rect 207980 9650 208000 9850
rect 204000 9640 208000 9650
rect 204140 9590 204360 9640
rect 204140 9520 204150 9590
rect 204350 9520 204360 9590
rect 204140 9480 204360 9520
rect 204140 9410 204150 9480
rect 204350 9410 204360 9480
rect 204140 9360 204360 9410
rect 204640 9590 204860 9640
rect 204640 9520 204650 9590
rect 204850 9520 204860 9590
rect 204640 9480 204860 9520
rect 204640 9410 204650 9480
rect 204850 9410 204860 9480
rect 204640 9360 204860 9410
rect 205140 9590 205360 9640
rect 205140 9520 205150 9590
rect 205350 9520 205360 9590
rect 205140 9480 205360 9520
rect 205140 9410 205150 9480
rect 205350 9410 205360 9480
rect 205140 9360 205360 9410
rect 205640 9590 205860 9640
rect 205640 9520 205650 9590
rect 205850 9520 205860 9590
rect 205640 9480 205860 9520
rect 205640 9410 205650 9480
rect 205850 9410 205860 9480
rect 205640 9360 205860 9410
rect 206140 9590 206360 9640
rect 206140 9520 206150 9590
rect 206350 9520 206360 9590
rect 206140 9480 206360 9520
rect 206140 9410 206150 9480
rect 206350 9410 206360 9480
rect 206140 9360 206360 9410
rect 206640 9590 206860 9640
rect 206640 9520 206650 9590
rect 206850 9520 206860 9590
rect 206640 9480 206860 9520
rect 206640 9410 206650 9480
rect 206850 9410 206860 9480
rect 206640 9360 206860 9410
rect 207140 9590 207360 9640
rect 207140 9520 207150 9590
rect 207350 9520 207360 9590
rect 207140 9480 207360 9520
rect 207140 9410 207150 9480
rect 207350 9410 207360 9480
rect 207140 9360 207360 9410
rect 207640 9590 207860 9640
rect 207640 9520 207650 9590
rect 207850 9520 207860 9590
rect 207640 9480 207860 9520
rect 207640 9410 207650 9480
rect 207850 9410 207860 9480
rect 207640 9360 207860 9410
rect 204000 9350 208000 9360
rect 204000 9150 204020 9350
rect 204090 9150 204410 9350
rect 204480 9150 204520 9350
rect 204590 9150 204910 9350
rect 204980 9150 205020 9350
rect 205090 9150 205410 9350
rect 205480 9150 205520 9350
rect 205590 9150 205910 9350
rect 205980 9150 206020 9350
rect 206090 9150 206410 9350
rect 206480 9150 206520 9350
rect 206590 9150 206910 9350
rect 206980 9150 207020 9350
rect 207090 9150 207410 9350
rect 207480 9150 207520 9350
rect 207590 9150 207910 9350
rect 207980 9150 208000 9350
rect 204000 9140 208000 9150
rect 204140 9090 204360 9140
rect 204140 9020 204150 9090
rect 204350 9020 204360 9090
rect 204140 8980 204360 9020
rect 204140 8910 204150 8980
rect 204350 8910 204360 8980
rect 204140 8860 204360 8910
rect 204640 9090 204860 9140
rect 204640 9020 204650 9090
rect 204850 9020 204860 9090
rect 204640 8980 204860 9020
rect 204640 8910 204650 8980
rect 204850 8910 204860 8980
rect 204640 8860 204860 8910
rect 205140 9090 205360 9140
rect 205140 9020 205150 9090
rect 205350 9020 205360 9090
rect 205140 8980 205360 9020
rect 205140 8910 205150 8980
rect 205350 8910 205360 8980
rect 205140 8860 205360 8910
rect 205640 9090 205860 9140
rect 205640 9020 205650 9090
rect 205850 9020 205860 9090
rect 205640 8980 205860 9020
rect 205640 8910 205650 8980
rect 205850 8910 205860 8980
rect 205640 8860 205860 8910
rect 206140 9090 206360 9140
rect 206140 9020 206150 9090
rect 206350 9020 206360 9090
rect 206140 8980 206360 9020
rect 206140 8910 206150 8980
rect 206350 8910 206360 8980
rect 206140 8860 206360 8910
rect 206640 9090 206860 9140
rect 206640 9020 206650 9090
rect 206850 9020 206860 9090
rect 206640 8980 206860 9020
rect 206640 8910 206650 8980
rect 206850 8910 206860 8980
rect 206640 8860 206860 8910
rect 207140 9090 207360 9140
rect 207140 9020 207150 9090
rect 207350 9020 207360 9090
rect 207140 8980 207360 9020
rect 207140 8910 207150 8980
rect 207350 8910 207360 8980
rect 207140 8860 207360 8910
rect 207640 9090 207860 9140
rect 207640 9020 207650 9090
rect 207850 9020 207860 9090
rect 207640 8980 207860 9020
rect 207640 8910 207650 8980
rect 207850 8910 207860 8980
rect 207640 8860 207860 8910
rect 204000 8850 208000 8860
rect 204000 8650 204020 8850
rect 204090 8650 204410 8850
rect 204480 8650 204520 8850
rect 204590 8650 204910 8850
rect 204980 8650 205020 8850
rect 205090 8650 205410 8850
rect 205480 8650 205520 8850
rect 205590 8650 205910 8850
rect 205980 8650 206020 8850
rect 206090 8650 206410 8850
rect 206480 8650 206520 8850
rect 206590 8650 206910 8850
rect 206980 8650 207020 8850
rect 207090 8650 207410 8850
rect 207480 8650 207520 8850
rect 207590 8650 207910 8850
rect 207980 8650 208000 8850
rect 204000 8640 208000 8650
rect 204140 8590 204360 8640
rect 204140 8520 204150 8590
rect 204350 8520 204360 8590
rect 204140 8480 204360 8520
rect 204140 8410 204150 8480
rect 204350 8410 204360 8480
rect 204140 8360 204360 8410
rect 204640 8590 204860 8640
rect 204640 8520 204650 8590
rect 204850 8520 204860 8590
rect 204640 8480 204860 8520
rect 204640 8410 204650 8480
rect 204850 8410 204860 8480
rect 204640 8360 204860 8410
rect 205140 8590 205360 8640
rect 205140 8520 205150 8590
rect 205350 8520 205360 8590
rect 205140 8480 205360 8520
rect 205140 8410 205150 8480
rect 205350 8410 205360 8480
rect 205140 8360 205360 8410
rect 205640 8590 205860 8640
rect 205640 8520 205650 8590
rect 205850 8520 205860 8590
rect 205640 8480 205860 8520
rect 205640 8410 205650 8480
rect 205850 8410 205860 8480
rect 205640 8360 205860 8410
rect 206140 8590 206360 8640
rect 206140 8520 206150 8590
rect 206350 8520 206360 8590
rect 206140 8480 206360 8520
rect 206140 8410 206150 8480
rect 206350 8410 206360 8480
rect 206140 8360 206360 8410
rect 206640 8590 206860 8640
rect 206640 8520 206650 8590
rect 206850 8520 206860 8590
rect 206640 8480 206860 8520
rect 206640 8410 206650 8480
rect 206850 8410 206860 8480
rect 206640 8360 206860 8410
rect 207140 8590 207360 8640
rect 207140 8520 207150 8590
rect 207350 8520 207360 8590
rect 207140 8480 207360 8520
rect 207140 8410 207150 8480
rect 207350 8410 207360 8480
rect 207140 8360 207360 8410
rect 207640 8590 207860 8640
rect 207640 8520 207650 8590
rect 207850 8520 207860 8590
rect 207640 8480 207860 8520
rect 207640 8410 207650 8480
rect 207850 8410 207860 8480
rect 207640 8360 207860 8410
rect 204000 8350 208000 8360
rect 204000 8150 204020 8350
rect 204090 8150 204410 8350
rect 204480 8150 204520 8350
rect 204590 8150 204910 8350
rect 204980 8150 205020 8350
rect 205090 8150 205410 8350
rect 205480 8150 205520 8350
rect 205590 8150 205910 8350
rect 205980 8150 206020 8350
rect 206090 8150 206410 8350
rect 206480 8150 206520 8350
rect 206590 8150 206910 8350
rect 206980 8150 207020 8350
rect 207090 8150 207410 8350
rect 207480 8150 207520 8350
rect 207590 8150 207910 8350
rect 207980 8150 208000 8350
rect 204000 8140 208000 8150
rect 204140 8090 204360 8140
rect 204140 8020 204150 8090
rect 204350 8020 204360 8090
rect 204140 7980 204360 8020
rect 204140 7910 204150 7980
rect 204350 7910 204360 7980
rect 204140 7860 204360 7910
rect 204640 8090 204860 8140
rect 204640 8020 204650 8090
rect 204850 8020 204860 8090
rect 204640 7980 204860 8020
rect 204640 7910 204650 7980
rect 204850 7910 204860 7980
rect 204640 7860 204860 7910
rect 205140 8090 205360 8140
rect 205140 8020 205150 8090
rect 205350 8020 205360 8090
rect 205140 7980 205360 8020
rect 205140 7910 205150 7980
rect 205350 7910 205360 7980
rect 205140 7860 205360 7910
rect 205640 8090 205860 8140
rect 205640 8020 205650 8090
rect 205850 8020 205860 8090
rect 205640 7980 205860 8020
rect 205640 7910 205650 7980
rect 205850 7910 205860 7980
rect 205640 7860 205860 7910
rect 206140 8090 206360 8140
rect 206140 8020 206150 8090
rect 206350 8020 206360 8090
rect 206140 7980 206360 8020
rect 206140 7910 206150 7980
rect 206350 7910 206360 7980
rect 206140 7860 206360 7910
rect 206640 8090 206860 8140
rect 206640 8020 206650 8090
rect 206850 8020 206860 8090
rect 206640 7980 206860 8020
rect 206640 7910 206650 7980
rect 206850 7910 206860 7980
rect 206640 7860 206860 7910
rect 207140 8090 207360 8140
rect 207140 8020 207150 8090
rect 207350 8020 207360 8090
rect 207140 7980 207360 8020
rect 207140 7910 207150 7980
rect 207350 7910 207360 7980
rect 207140 7860 207360 7910
rect 207640 8090 207860 8140
rect 207640 8020 207650 8090
rect 207850 8020 207860 8090
rect 207640 7980 207860 8020
rect 207640 7910 207650 7980
rect 207850 7910 207860 7980
rect 207640 7860 207860 7910
rect 204000 7850 208000 7860
rect 204000 7650 204020 7850
rect 204090 7650 204410 7850
rect 204480 7650 204520 7850
rect 204590 7650 204910 7850
rect 204980 7650 205020 7850
rect 205090 7650 205410 7850
rect 205480 7650 205520 7850
rect 205590 7650 205910 7850
rect 205980 7650 206020 7850
rect 206090 7650 206410 7850
rect 206480 7650 206520 7850
rect 206590 7650 206910 7850
rect 206980 7650 207020 7850
rect 207090 7650 207410 7850
rect 207480 7650 207520 7850
rect 207590 7650 207910 7850
rect 207980 7650 208000 7850
rect 204000 7640 208000 7650
rect 204140 7590 204360 7640
rect 204140 7520 204150 7590
rect 204350 7520 204360 7590
rect 204140 7480 204360 7520
rect 204140 7410 204150 7480
rect 204350 7410 204360 7480
rect 204140 7360 204360 7410
rect 204640 7590 204860 7640
rect 204640 7520 204650 7590
rect 204850 7520 204860 7590
rect 204640 7480 204860 7520
rect 204640 7410 204650 7480
rect 204850 7410 204860 7480
rect 204640 7360 204860 7410
rect 205140 7590 205360 7640
rect 205140 7520 205150 7590
rect 205350 7520 205360 7590
rect 205140 7480 205360 7520
rect 205140 7410 205150 7480
rect 205350 7410 205360 7480
rect 205140 7360 205360 7410
rect 205640 7590 205860 7640
rect 205640 7520 205650 7590
rect 205850 7520 205860 7590
rect 205640 7480 205860 7520
rect 205640 7410 205650 7480
rect 205850 7410 205860 7480
rect 205640 7360 205860 7410
rect 206140 7590 206360 7640
rect 206140 7520 206150 7590
rect 206350 7520 206360 7590
rect 206140 7480 206360 7520
rect 206140 7410 206150 7480
rect 206350 7410 206360 7480
rect 206140 7360 206360 7410
rect 206640 7590 206860 7640
rect 206640 7520 206650 7590
rect 206850 7520 206860 7590
rect 206640 7480 206860 7520
rect 206640 7410 206650 7480
rect 206850 7410 206860 7480
rect 206640 7360 206860 7410
rect 207140 7590 207360 7640
rect 207140 7520 207150 7590
rect 207350 7520 207360 7590
rect 207140 7480 207360 7520
rect 207140 7410 207150 7480
rect 207350 7410 207360 7480
rect 207140 7360 207360 7410
rect 207640 7590 207860 7640
rect 207640 7520 207650 7590
rect 207850 7520 207860 7590
rect 207640 7480 207860 7520
rect 207640 7410 207650 7480
rect 207850 7410 207860 7480
rect 207640 7360 207860 7410
rect 204000 7350 208000 7360
rect 204000 7150 204020 7350
rect 204090 7150 204410 7350
rect 204480 7150 204520 7350
rect 204590 7150 204910 7350
rect 204980 7150 205020 7350
rect 205090 7150 205410 7350
rect 205480 7150 205520 7350
rect 205590 7150 205910 7350
rect 205980 7150 206020 7350
rect 206090 7150 206410 7350
rect 206480 7150 206520 7350
rect 206590 7150 206910 7350
rect 206980 7150 207020 7350
rect 207090 7150 207410 7350
rect 207480 7150 207520 7350
rect 207590 7150 207910 7350
rect 207980 7150 208000 7350
rect 204000 7140 208000 7150
rect 204140 7090 204360 7140
rect 204140 7020 204150 7090
rect 204350 7020 204360 7090
rect 204140 6980 204360 7020
rect 204140 6910 204150 6980
rect 204350 6910 204360 6980
rect 204140 6860 204360 6910
rect 204640 7090 204860 7140
rect 204640 7020 204650 7090
rect 204850 7020 204860 7090
rect 204640 6980 204860 7020
rect 204640 6910 204650 6980
rect 204850 6910 204860 6980
rect 204640 6860 204860 6910
rect 205140 7090 205360 7140
rect 205140 7020 205150 7090
rect 205350 7020 205360 7090
rect 205140 6980 205360 7020
rect 205140 6910 205150 6980
rect 205350 6910 205360 6980
rect 205140 6860 205360 6910
rect 205640 7090 205860 7140
rect 205640 7020 205650 7090
rect 205850 7020 205860 7090
rect 205640 6980 205860 7020
rect 205640 6910 205650 6980
rect 205850 6910 205860 6980
rect 205640 6860 205860 6910
rect 206140 7090 206360 7140
rect 206140 7020 206150 7090
rect 206350 7020 206360 7090
rect 206140 6980 206360 7020
rect 206140 6910 206150 6980
rect 206350 6910 206360 6980
rect 206140 6860 206360 6910
rect 206640 7090 206860 7140
rect 206640 7020 206650 7090
rect 206850 7020 206860 7090
rect 206640 6980 206860 7020
rect 206640 6910 206650 6980
rect 206850 6910 206860 6980
rect 206640 6860 206860 6910
rect 207140 7090 207360 7140
rect 207140 7020 207150 7090
rect 207350 7020 207360 7090
rect 207140 6980 207360 7020
rect 207140 6910 207150 6980
rect 207350 6910 207360 6980
rect 207140 6860 207360 6910
rect 207640 7090 207860 7140
rect 207640 7020 207650 7090
rect 207850 7020 207860 7090
rect 207640 6980 207860 7020
rect 207640 6910 207650 6980
rect 207850 6910 207860 6980
rect 207640 6860 207860 6910
rect 204000 6850 208000 6860
rect 204000 6650 204020 6850
rect 204090 6650 204410 6850
rect 204480 6650 204520 6850
rect 204590 6650 204910 6850
rect 204980 6650 205020 6850
rect 205090 6650 205410 6850
rect 205480 6650 205520 6850
rect 205590 6650 205910 6850
rect 205980 6650 206020 6850
rect 206090 6650 206410 6850
rect 206480 6650 206520 6850
rect 206590 6650 206910 6850
rect 206980 6650 207020 6850
rect 207090 6650 207410 6850
rect 207480 6650 207520 6850
rect 207590 6650 207910 6850
rect 207980 6650 208000 6850
rect 204000 6640 208000 6650
rect 204140 6590 204360 6640
rect 204140 6520 204150 6590
rect 204350 6520 204360 6590
rect 204140 6480 204360 6520
rect 204140 6410 204150 6480
rect 204350 6410 204360 6480
rect 204140 6360 204360 6410
rect 204640 6590 204860 6640
rect 204640 6520 204650 6590
rect 204850 6520 204860 6590
rect 204640 6480 204860 6520
rect 204640 6410 204650 6480
rect 204850 6410 204860 6480
rect 204640 6360 204860 6410
rect 205140 6590 205360 6640
rect 205140 6520 205150 6590
rect 205350 6520 205360 6590
rect 205140 6480 205360 6520
rect 205140 6410 205150 6480
rect 205350 6410 205360 6480
rect 205140 6360 205360 6410
rect 205640 6590 205860 6640
rect 205640 6520 205650 6590
rect 205850 6520 205860 6590
rect 205640 6480 205860 6520
rect 205640 6410 205650 6480
rect 205850 6410 205860 6480
rect 205640 6360 205860 6410
rect 206140 6590 206360 6640
rect 206140 6520 206150 6590
rect 206350 6520 206360 6590
rect 206140 6480 206360 6520
rect 206140 6410 206150 6480
rect 206350 6410 206360 6480
rect 206140 6360 206360 6410
rect 206640 6590 206860 6640
rect 206640 6520 206650 6590
rect 206850 6520 206860 6590
rect 206640 6480 206860 6520
rect 206640 6410 206650 6480
rect 206850 6410 206860 6480
rect 206640 6360 206860 6410
rect 207140 6590 207360 6640
rect 207140 6520 207150 6590
rect 207350 6520 207360 6590
rect 207140 6480 207360 6520
rect 207140 6410 207150 6480
rect 207350 6410 207360 6480
rect 207140 6360 207360 6410
rect 207640 6590 207860 6640
rect 207640 6520 207650 6590
rect 207850 6520 207860 6590
rect 207640 6480 207860 6520
rect 207640 6410 207650 6480
rect 207850 6410 207860 6480
rect 207640 6360 207860 6410
rect 204000 6350 208000 6360
rect 204000 6150 204020 6350
rect 204090 6150 204410 6350
rect 204480 6150 204520 6350
rect 204590 6150 204910 6350
rect 204980 6150 205020 6350
rect 205090 6150 205410 6350
rect 205480 6150 205520 6350
rect 205590 6150 205910 6350
rect 205980 6150 206020 6350
rect 206090 6150 206410 6350
rect 206480 6150 206520 6350
rect 206590 6150 206910 6350
rect 206980 6150 207020 6350
rect 207090 6150 207410 6350
rect 207480 6150 207520 6350
rect 207590 6150 207910 6350
rect 207980 6150 208000 6350
rect 204000 6140 208000 6150
rect 204140 6090 204360 6140
rect 204140 6020 204150 6090
rect 204350 6020 204360 6090
rect 198140 5980 198360 6000
rect 198140 5910 198150 5980
rect 198350 5910 198360 5980
rect 198140 5860 198360 5910
rect 198640 5980 198860 6000
rect 198640 5910 198650 5980
rect 198850 5910 198860 5980
rect 198640 5860 198860 5910
rect 199140 5980 199360 6000
rect 199140 5910 199150 5980
rect 199350 5910 199360 5980
rect 199140 5860 199360 5910
rect 199640 5980 199860 6000
rect 199640 5910 199650 5980
rect 199850 5910 199860 5980
rect 199640 5860 199860 5910
rect 200140 5980 200360 6000
rect 200140 5910 200150 5980
rect 200350 5910 200360 5980
rect 200140 5860 200360 5910
rect 200640 5980 200860 6000
rect 200640 5910 200650 5980
rect 200850 5910 200860 5980
rect 200640 5860 200860 5910
rect 201140 5980 201360 6000
rect 201140 5910 201150 5980
rect 201350 5910 201360 5980
rect 201140 5860 201360 5910
rect 201640 5980 201860 6000
rect 201640 5910 201650 5980
rect 201850 5910 201860 5980
rect 201640 5860 201860 5910
rect 202140 5980 202360 6000
rect 202140 5910 202150 5980
rect 202350 5910 202360 5980
rect 202140 5860 202360 5910
rect 202640 5980 202860 6000
rect 202640 5910 202650 5980
rect 202850 5910 202860 5980
rect 202640 5860 202860 5910
rect 203140 5980 203360 6000
rect 203140 5910 203150 5980
rect 203350 5910 203360 5980
rect 203140 5860 203360 5910
rect 203640 5980 203860 6000
rect 203640 5910 203650 5980
rect 203850 5910 203860 5980
rect 203640 5860 203860 5910
rect 204140 5980 204360 6020
rect 204140 5910 204150 5980
rect 204350 5910 204360 5980
rect 204140 5860 204360 5910
rect 204640 6090 204860 6140
rect 204640 6020 204650 6090
rect 204850 6020 204860 6090
rect 204640 5980 204860 6020
rect 204640 5910 204650 5980
rect 204850 5910 204860 5980
rect 204640 5860 204860 5910
rect 205140 6090 205360 6140
rect 205140 6020 205150 6090
rect 205350 6020 205360 6090
rect 205140 5980 205360 6020
rect 205140 5910 205150 5980
rect 205350 5910 205360 5980
rect 205140 5860 205360 5910
rect 205640 6090 205860 6140
rect 205640 6020 205650 6090
rect 205850 6020 205860 6090
rect 205640 5980 205860 6020
rect 205640 5910 205650 5980
rect 205850 5910 205860 5980
rect 205640 5860 205860 5910
rect 206140 6090 206360 6140
rect 206140 6020 206150 6090
rect 206350 6020 206360 6090
rect 206140 5980 206360 6020
rect 206140 5910 206150 5980
rect 206350 5910 206360 5980
rect 206140 5860 206360 5910
rect 206640 6090 206860 6140
rect 206640 6020 206650 6090
rect 206850 6020 206860 6090
rect 206640 5980 206860 6020
rect 206640 5910 206650 5980
rect 206850 5910 206860 5980
rect 206640 5860 206860 5910
rect 207140 6090 207360 6140
rect 207140 6020 207150 6090
rect 207350 6020 207360 6090
rect 207140 5980 207360 6020
rect 207140 5910 207150 5980
rect 207350 5910 207360 5980
rect 207140 5860 207360 5910
rect 207640 6090 207860 6140
rect 207640 6020 207650 6090
rect 207850 6020 207860 6090
rect 207640 5980 207860 6020
rect 207640 5910 207650 5980
rect 207850 5910 207860 5980
rect 207640 5860 207860 5910
rect 198000 5850 208000 5860
rect 198000 5650 198020 5850
rect 198090 5650 198410 5850
rect 198480 5650 198520 5850
rect 198590 5650 198910 5850
rect 198980 5650 199020 5850
rect 199090 5650 199410 5850
rect 199480 5650 199520 5850
rect 199590 5650 199910 5850
rect 199980 5650 200020 5850
rect 200090 5650 200410 5850
rect 200480 5650 200520 5850
rect 200590 5650 200910 5850
rect 200980 5650 201020 5850
rect 201090 5650 201410 5850
rect 201480 5650 201520 5850
rect 201590 5650 201910 5850
rect 201980 5650 202020 5850
rect 202090 5650 202410 5850
rect 202480 5650 202520 5850
rect 202590 5650 202910 5850
rect 202980 5650 203020 5850
rect 203090 5650 203410 5850
rect 203480 5650 203520 5850
rect 203590 5650 203910 5850
rect 203980 5650 204020 5850
rect 204090 5650 204410 5850
rect 204480 5650 204520 5850
rect 204590 5650 204910 5850
rect 204980 5650 205020 5850
rect 205090 5650 205410 5850
rect 205480 5650 205520 5850
rect 205590 5650 205910 5850
rect 205980 5650 206020 5850
rect 206090 5650 206410 5850
rect 206480 5650 206520 5850
rect 206590 5650 206910 5850
rect 206980 5650 207020 5850
rect 207090 5650 207410 5850
rect 207480 5650 207520 5850
rect 207590 5650 207910 5850
rect 207980 5650 208000 5850
rect 198000 5640 208000 5650
rect 198140 5590 198360 5640
rect 198140 5520 198150 5590
rect 198350 5520 198360 5590
rect 198140 5480 198360 5520
rect 198140 5410 198150 5480
rect 198350 5410 198360 5480
rect 198140 5360 198360 5410
rect 198640 5590 198860 5640
rect 198640 5520 198650 5590
rect 198850 5520 198860 5590
rect 198640 5480 198860 5520
rect 198640 5410 198650 5480
rect 198850 5410 198860 5480
rect 198640 5360 198860 5410
rect 199140 5590 199360 5640
rect 199140 5520 199150 5590
rect 199350 5520 199360 5590
rect 199140 5480 199360 5520
rect 199140 5410 199150 5480
rect 199350 5410 199360 5480
rect 199140 5360 199360 5410
rect 199640 5590 199860 5640
rect 199640 5520 199650 5590
rect 199850 5520 199860 5590
rect 199640 5480 199860 5520
rect 199640 5410 199650 5480
rect 199850 5410 199860 5480
rect 199640 5360 199860 5410
rect 200140 5590 200360 5640
rect 200140 5520 200150 5590
rect 200350 5520 200360 5590
rect 200140 5480 200360 5520
rect 200140 5410 200150 5480
rect 200350 5410 200360 5480
rect 200140 5360 200360 5410
rect 200640 5590 200860 5640
rect 200640 5520 200650 5590
rect 200850 5520 200860 5590
rect 200640 5480 200860 5520
rect 200640 5410 200650 5480
rect 200850 5410 200860 5480
rect 200640 5360 200860 5410
rect 201140 5590 201360 5640
rect 201140 5520 201150 5590
rect 201350 5520 201360 5590
rect 201140 5480 201360 5520
rect 201140 5410 201150 5480
rect 201350 5410 201360 5480
rect 201140 5360 201360 5410
rect 201640 5590 201860 5640
rect 201640 5520 201650 5590
rect 201850 5520 201860 5590
rect 201640 5480 201860 5520
rect 201640 5410 201650 5480
rect 201850 5410 201860 5480
rect 201640 5360 201860 5410
rect 202140 5590 202360 5640
rect 202140 5520 202150 5590
rect 202350 5520 202360 5590
rect 202140 5480 202360 5520
rect 202140 5410 202150 5480
rect 202350 5410 202360 5480
rect 202140 5360 202360 5410
rect 202640 5590 202860 5640
rect 202640 5520 202650 5590
rect 202850 5520 202860 5590
rect 202640 5480 202860 5520
rect 202640 5410 202650 5480
rect 202850 5410 202860 5480
rect 202640 5360 202860 5410
rect 203140 5590 203360 5640
rect 203140 5520 203150 5590
rect 203350 5520 203360 5590
rect 203140 5480 203360 5520
rect 203140 5410 203150 5480
rect 203350 5410 203360 5480
rect 203140 5360 203360 5410
rect 203640 5590 203860 5640
rect 203640 5520 203650 5590
rect 203850 5520 203860 5590
rect 203640 5480 203860 5520
rect 203640 5410 203650 5480
rect 203850 5410 203860 5480
rect 203640 5360 203860 5410
rect 204140 5590 204360 5640
rect 204140 5520 204150 5590
rect 204350 5520 204360 5590
rect 204140 5480 204360 5520
rect 204140 5410 204150 5480
rect 204350 5410 204360 5480
rect 204140 5360 204360 5410
rect 204640 5590 204860 5640
rect 204640 5520 204650 5590
rect 204850 5520 204860 5590
rect 204640 5480 204860 5520
rect 204640 5410 204650 5480
rect 204850 5410 204860 5480
rect 204640 5360 204860 5410
rect 205140 5590 205360 5640
rect 205140 5520 205150 5590
rect 205350 5520 205360 5590
rect 205140 5480 205360 5520
rect 205140 5410 205150 5480
rect 205350 5410 205360 5480
rect 205140 5360 205360 5410
rect 205640 5590 205860 5640
rect 205640 5520 205650 5590
rect 205850 5520 205860 5590
rect 205640 5480 205860 5520
rect 205640 5410 205650 5480
rect 205850 5410 205860 5480
rect 205640 5360 205860 5410
rect 206140 5590 206360 5640
rect 206140 5520 206150 5590
rect 206350 5520 206360 5590
rect 206140 5480 206360 5520
rect 206140 5410 206150 5480
rect 206350 5410 206360 5480
rect 206140 5360 206360 5410
rect 206640 5590 206860 5640
rect 206640 5520 206650 5590
rect 206850 5520 206860 5590
rect 206640 5480 206860 5520
rect 206640 5410 206650 5480
rect 206850 5410 206860 5480
rect 206640 5360 206860 5410
rect 207140 5590 207360 5640
rect 207140 5520 207150 5590
rect 207350 5520 207360 5590
rect 207140 5480 207360 5520
rect 207140 5410 207150 5480
rect 207350 5410 207360 5480
rect 207140 5360 207360 5410
rect 207640 5590 207860 5640
rect 207640 5520 207650 5590
rect 207850 5520 207860 5590
rect 207640 5480 207860 5520
rect 207640 5410 207650 5480
rect 207850 5410 207860 5480
rect 207640 5360 207860 5410
rect 198000 5350 208000 5360
rect 198000 5150 198020 5350
rect 198090 5150 198410 5350
rect 198480 5150 198520 5350
rect 198590 5150 198910 5350
rect 198980 5150 199020 5350
rect 199090 5150 199410 5350
rect 199480 5150 199520 5350
rect 199590 5150 199910 5350
rect 199980 5150 200020 5350
rect 200090 5150 200410 5350
rect 200480 5150 200520 5350
rect 200590 5150 200910 5350
rect 200980 5150 201020 5350
rect 201090 5150 201410 5350
rect 201480 5150 201520 5350
rect 201590 5150 201910 5350
rect 201980 5150 202020 5350
rect 202090 5150 202410 5350
rect 202480 5150 202520 5350
rect 202590 5150 202910 5350
rect 202980 5150 203020 5350
rect 203090 5150 203410 5350
rect 203480 5150 203520 5350
rect 203590 5150 203910 5350
rect 203980 5150 204020 5350
rect 204090 5150 204410 5350
rect 204480 5150 204520 5350
rect 204590 5150 204910 5350
rect 204980 5150 205020 5350
rect 205090 5150 205410 5350
rect 205480 5150 205520 5350
rect 205590 5150 205910 5350
rect 205980 5150 206020 5350
rect 206090 5150 206410 5350
rect 206480 5150 206520 5350
rect 206590 5150 206910 5350
rect 206980 5150 207020 5350
rect 207090 5150 207410 5350
rect 207480 5150 207520 5350
rect 207590 5150 207910 5350
rect 207980 5150 208000 5350
rect 198000 5140 208000 5150
rect 198140 5090 198360 5140
rect 198140 5020 198150 5090
rect 198350 5020 198360 5090
rect 198140 4980 198360 5020
rect 198140 4910 198150 4980
rect 198350 4910 198360 4980
rect 198140 4860 198360 4910
rect 198640 5090 198860 5140
rect 198640 5020 198650 5090
rect 198850 5020 198860 5090
rect 198640 4980 198860 5020
rect 198640 4910 198650 4980
rect 198850 4910 198860 4980
rect 198640 4860 198860 4910
rect 199140 5090 199360 5140
rect 199140 5020 199150 5090
rect 199350 5020 199360 5090
rect 199140 4980 199360 5020
rect 199140 4910 199150 4980
rect 199350 4910 199360 4980
rect 199140 4860 199360 4910
rect 199640 5090 199860 5140
rect 199640 5020 199650 5090
rect 199850 5020 199860 5090
rect 199640 4980 199860 5020
rect 199640 4910 199650 4980
rect 199850 4910 199860 4980
rect 199640 4860 199860 4910
rect 200140 5090 200360 5140
rect 200140 5020 200150 5090
rect 200350 5020 200360 5090
rect 200140 4980 200360 5020
rect 200140 4910 200150 4980
rect 200350 4910 200360 4980
rect 200140 4860 200360 4910
rect 200640 5090 200860 5140
rect 200640 5020 200650 5090
rect 200850 5020 200860 5090
rect 200640 4980 200860 5020
rect 200640 4910 200650 4980
rect 200850 4910 200860 4980
rect 200640 4860 200860 4910
rect 201140 5090 201360 5140
rect 201140 5020 201150 5090
rect 201350 5020 201360 5090
rect 201140 4980 201360 5020
rect 201140 4910 201150 4980
rect 201350 4910 201360 4980
rect 201140 4860 201360 4910
rect 201640 5090 201860 5140
rect 201640 5020 201650 5090
rect 201850 5020 201860 5090
rect 201640 4980 201860 5020
rect 201640 4910 201650 4980
rect 201850 4910 201860 4980
rect 201640 4860 201860 4910
rect 202140 5090 202360 5140
rect 202140 5020 202150 5090
rect 202350 5020 202360 5090
rect 202140 4980 202360 5020
rect 202140 4910 202150 4980
rect 202350 4910 202360 4980
rect 202140 4860 202360 4910
rect 202640 5090 202860 5140
rect 202640 5020 202650 5090
rect 202850 5020 202860 5090
rect 202640 4980 202860 5020
rect 202640 4910 202650 4980
rect 202850 4910 202860 4980
rect 202640 4860 202860 4910
rect 203140 5090 203360 5140
rect 203140 5020 203150 5090
rect 203350 5020 203360 5090
rect 203140 4980 203360 5020
rect 203140 4910 203150 4980
rect 203350 4910 203360 4980
rect 203140 4860 203360 4910
rect 203640 5090 203860 5140
rect 203640 5020 203650 5090
rect 203850 5020 203860 5090
rect 203640 4980 203860 5020
rect 203640 4910 203650 4980
rect 203850 4910 203860 4980
rect 203640 4860 203860 4910
rect 204140 5090 204360 5140
rect 204140 5020 204150 5090
rect 204350 5020 204360 5090
rect 204140 4980 204360 5020
rect 204140 4910 204150 4980
rect 204350 4910 204360 4980
rect 204140 4860 204360 4910
rect 204640 5090 204860 5140
rect 204640 5020 204650 5090
rect 204850 5020 204860 5090
rect 204640 4980 204860 5020
rect 204640 4910 204650 4980
rect 204850 4910 204860 4980
rect 204640 4860 204860 4910
rect 205140 5090 205360 5140
rect 205140 5020 205150 5090
rect 205350 5020 205360 5090
rect 205140 4980 205360 5020
rect 205140 4910 205150 4980
rect 205350 4910 205360 4980
rect 205140 4860 205360 4910
rect 205640 5090 205860 5140
rect 205640 5020 205650 5090
rect 205850 5020 205860 5090
rect 205640 4980 205860 5020
rect 205640 4910 205650 4980
rect 205850 4910 205860 4980
rect 205640 4860 205860 4910
rect 206140 5090 206360 5140
rect 206140 5020 206150 5090
rect 206350 5020 206360 5090
rect 206140 4980 206360 5020
rect 206140 4910 206150 4980
rect 206350 4910 206360 4980
rect 206140 4860 206360 4910
rect 206640 5090 206860 5140
rect 206640 5020 206650 5090
rect 206850 5020 206860 5090
rect 206640 4980 206860 5020
rect 206640 4910 206650 4980
rect 206850 4910 206860 4980
rect 206640 4860 206860 4910
rect 207140 5090 207360 5140
rect 207140 5020 207150 5090
rect 207350 5020 207360 5090
rect 207140 4980 207360 5020
rect 207140 4910 207150 4980
rect 207350 4910 207360 4980
rect 207140 4860 207360 4910
rect 207640 5090 207860 5140
rect 207640 5020 207650 5090
rect 207850 5020 207860 5090
rect 207640 4980 207860 5020
rect 207640 4910 207650 4980
rect 207850 4910 207860 4980
rect 207640 4860 207860 4910
rect 198000 4850 208000 4860
rect 198000 4650 198020 4850
rect 198090 4650 198410 4850
rect 198480 4650 198520 4850
rect 198590 4650 198910 4850
rect 198980 4650 199020 4850
rect 199090 4650 199410 4850
rect 199480 4650 199520 4850
rect 199590 4650 199910 4850
rect 199980 4650 200020 4850
rect 200090 4650 200410 4850
rect 200480 4650 200520 4850
rect 200590 4650 200910 4850
rect 200980 4650 201020 4850
rect 201090 4650 201410 4850
rect 201480 4650 201520 4850
rect 201590 4650 201910 4850
rect 201980 4650 202020 4850
rect 202090 4650 202410 4850
rect 202480 4650 202520 4850
rect 202590 4650 202910 4850
rect 202980 4650 203020 4850
rect 203090 4650 203410 4850
rect 203480 4650 203520 4850
rect 203590 4650 203910 4850
rect 203980 4650 204020 4850
rect 204090 4650 204410 4850
rect 204480 4650 204520 4850
rect 204590 4650 204910 4850
rect 204980 4650 205020 4850
rect 205090 4650 205410 4850
rect 205480 4650 205520 4850
rect 205590 4650 205910 4850
rect 205980 4650 206020 4850
rect 206090 4650 206410 4850
rect 206480 4650 206520 4850
rect 206590 4650 206910 4850
rect 206980 4650 207020 4850
rect 207090 4650 207410 4850
rect 207480 4650 207520 4850
rect 207590 4650 207910 4850
rect 207980 4650 208000 4850
rect 198000 4640 208000 4650
rect 198140 4590 198360 4640
rect 198140 4520 198150 4590
rect 198350 4520 198360 4590
rect 198140 4480 198360 4520
rect 198140 4410 198150 4480
rect 198350 4410 198360 4480
rect 198140 4360 198360 4410
rect 198640 4590 198860 4640
rect 198640 4520 198650 4590
rect 198850 4520 198860 4590
rect 198640 4480 198860 4520
rect 198640 4410 198650 4480
rect 198850 4410 198860 4480
rect 198640 4360 198860 4410
rect 199140 4590 199360 4640
rect 199140 4520 199150 4590
rect 199350 4520 199360 4590
rect 199140 4480 199360 4520
rect 199140 4410 199150 4480
rect 199350 4410 199360 4480
rect 199140 4360 199360 4410
rect 199640 4590 199860 4640
rect 199640 4520 199650 4590
rect 199850 4520 199860 4590
rect 199640 4480 199860 4520
rect 199640 4410 199650 4480
rect 199850 4410 199860 4480
rect 199640 4360 199860 4410
rect 200140 4590 200360 4640
rect 200140 4520 200150 4590
rect 200350 4520 200360 4590
rect 200140 4480 200360 4520
rect 200140 4410 200150 4480
rect 200350 4410 200360 4480
rect 200140 4360 200360 4410
rect 200640 4590 200860 4640
rect 200640 4520 200650 4590
rect 200850 4520 200860 4590
rect 200640 4480 200860 4520
rect 200640 4410 200650 4480
rect 200850 4410 200860 4480
rect 200640 4360 200860 4410
rect 201140 4590 201360 4640
rect 201140 4520 201150 4590
rect 201350 4520 201360 4590
rect 201140 4480 201360 4520
rect 201140 4410 201150 4480
rect 201350 4410 201360 4480
rect 201140 4360 201360 4410
rect 201640 4590 201860 4640
rect 201640 4520 201650 4590
rect 201850 4520 201860 4590
rect 201640 4480 201860 4520
rect 201640 4410 201650 4480
rect 201850 4410 201860 4480
rect 201640 4360 201860 4410
rect 202140 4590 202360 4640
rect 202140 4520 202150 4590
rect 202350 4520 202360 4590
rect 202140 4480 202360 4520
rect 202140 4410 202150 4480
rect 202350 4410 202360 4480
rect 202140 4360 202360 4410
rect 202640 4590 202860 4640
rect 202640 4520 202650 4590
rect 202850 4520 202860 4590
rect 202640 4480 202860 4520
rect 202640 4410 202650 4480
rect 202850 4410 202860 4480
rect 202640 4360 202860 4410
rect 203140 4590 203360 4640
rect 203140 4520 203150 4590
rect 203350 4520 203360 4590
rect 203140 4480 203360 4520
rect 203140 4410 203150 4480
rect 203350 4410 203360 4480
rect 203140 4360 203360 4410
rect 203640 4590 203860 4640
rect 203640 4520 203650 4590
rect 203850 4520 203860 4590
rect 203640 4480 203860 4520
rect 203640 4410 203650 4480
rect 203850 4410 203860 4480
rect 203640 4360 203860 4410
rect 204140 4590 204360 4640
rect 204140 4520 204150 4590
rect 204350 4520 204360 4590
rect 204140 4480 204360 4520
rect 204140 4410 204150 4480
rect 204350 4410 204360 4480
rect 204140 4360 204360 4410
rect 204640 4590 204860 4640
rect 204640 4520 204650 4590
rect 204850 4520 204860 4590
rect 204640 4480 204860 4520
rect 204640 4410 204650 4480
rect 204850 4410 204860 4480
rect 204640 4360 204860 4410
rect 205140 4590 205360 4640
rect 205140 4520 205150 4590
rect 205350 4520 205360 4590
rect 205140 4480 205360 4520
rect 205140 4410 205150 4480
rect 205350 4410 205360 4480
rect 205140 4360 205360 4410
rect 205640 4590 205860 4640
rect 205640 4520 205650 4590
rect 205850 4520 205860 4590
rect 205640 4480 205860 4520
rect 205640 4410 205650 4480
rect 205850 4410 205860 4480
rect 205640 4360 205860 4410
rect 206140 4590 206360 4640
rect 206140 4520 206150 4590
rect 206350 4520 206360 4590
rect 206140 4480 206360 4520
rect 206140 4410 206150 4480
rect 206350 4410 206360 4480
rect 206140 4360 206360 4410
rect 206640 4590 206860 4640
rect 206640 4520 206650 4590
rect 206850 4520 206860 4590
rect 206640 4480 206860 4520
rect 206640 4410 206650 4480
rect 206850 4410 206860 4480
rect 206640 4360 206860 4410
rect 207140 4590 207360 4640
rect 207140 4520 207150 4590
rect 207350 4520 207360 4590
rect 207140 4480 207360 4520
rect 207140 4410 207150 4480
rect 207350 4410 207360 4480
rect 207140 4360 207360 4410
rect 207640 4590 207860 4640
rect 207640 4520 207650 4590
rect 207850 4520 207860 4590
rect 207640 4480 207860 4520
rect 207640 4410 207650 4480
rect 207850 4410 207860 4480
rect 207640 4360 207860 4410
rect 198000 4350 208000 4360
rect 198000 4150 198020 4350
rect 198090 4150 198410 4350
rect 198480 4150 198520 4350
rect 198590 4150 198910 4350
rect 198980 4150 199020 4350
rect 199090 4150 199410 4350
rect 199480 4150 199520 4350
rect 199590 4150 199910 4350
rect 199980 4150 200020 4350
rect 200090 4150 200410 4350
rect 200480 4150 200520 4350
rect 200590 4150 200910 4350
rect 200980 4150 201020 4350
rect 201090 4150 201410 4350
rect 201480 4150 201520 4350
rect 201590 4150 201910 4350
rect 201980 4150 202020 4350
rect 202090 4150 202410 4350
rect 202480 4150 202520 4350
rect 202590 4150 202910 4350
rect 202980 4150 203020 4350
rect 203090 4150 203410 4350
rect 203480 4150 203520 4350
rect 203590 4150 203910 4350
rect 203980 4150 204020 4350
rect 204090 4150 204410 4350
rect 204480 4150 204520 4350
rect 204590 4150 204910 4350
rect 204980 4150 205020 4350
rect 205090 4150 205410 4350
rect 205480 4150 205520 4350
rect 205590 4150 205910 4350
rect 205980 4150 206020 4350
rect 206090 4150 206410 4350
rect 206480 4150 206520 4350
rect 206590 4150 206910 4350
rect 206980 4150 207020 4350
rect 207090 4150 207410 4350
rect 207480 4150 207520 4350
rect 207590 4150 207910 4350
rect 207980 4150 208000 4350
rect 198000 4140 208000 4150
rect 198140 4090 198360 4140
rect 198140 4020 198150 4090
rect 198350 4020 198360 4090
rect 198140 3980 198360 4020
rect 198140 3910 198150 3980
rect 198350 3910 198360 3980
rect 198140 3860 198360 3910
rect 198640 4090 198860 4140
rect 198640 4020 198650 4090
rect 198850 4020 198860 4090
rect 198640 3980 198860 4020
rect 198640 3910 198650 3980
rect 198850 3910 198860 3980
rect 198640 3860 198860 3910
rect 199140 4090 199360 4140
rect 199140 4020 199150 4090
rect 199350 4020 199360 4090
rect 199140 3980 199360 4020
rect 199140 3910 199150 3980
rect 199350 3910 199360 3980
rect 199140 3860 199360 3910
rect 199640 4090 199860 4140
rect 199640 4020 199650 4090
rect 199850 4020 199860 4090
rect 199640 3980 199860 4020
rect 199640 3910 199650 3980
rect 199850 3910 199860 3980
rect 199640 3860 199860 3910
rect 200140 4090 200360 4140
rect 200140 4020 200150 4090
rect 200350 4020 200360 4090
rect 200140 3980 200360 4020
rect 200140 3910 200150 3980
rect 200350 3910 200360 3980
rect 200140 3860 200360 3910
rect 200640 4090 200860 4140
rect 200640 4020 200650 4090
rect 200850 4020 200860 4090
rect 200640 3980 200860 4020
rect 200640 3910 200650 3980
rect 200850 3910 200860 3980
rect 200640 3860 200860 3910
rect 201140 4090 201360 4140
rect 201140 4020 201150 4090
rect 201350 4020 201360 4090
rect 201140 3980 201360 4020
rect 201140 3910 201150 3980
rect 201350 3910 201360 3980
rect 201140 3860 201360 3910
rect 201640 4090 201860 4140
rect 201640 4020 201650 4090
rect 201850 4020 201860 4090
rect 201640 3980 201860 4020
rect 201640 3910 201650 3980
rect 201850 3910 201860 3980
rect 201640 3860 201860 3910
rect 202140 4090 202360 4140
rect 202140 4020 202150 4090
rect 202350 4020 202360 4090
rect 202140 3980 202360 4020
rect 202140 3910 202150 3980
rect 202350 3910 202360 3980
rect 202140 3860 202360 3910
rect 202640 4090 202860 4140
rect 202640 4020 202650 4090
rect 202850 4020 202860 4090
rect 202640 3980 202860 4020
rect 202640 3910 202650 3980
rect 202850 3910 202860 3980
rect 202640 3860 202860 3910
rect 203140 4090 203360 4140
rect 203140 4020 203150 4090
rect 203350 4020 203360 4090
rect 203140 3980 203360 4020
rect 203140 3910 203150 3980
rect 203350 3910 203360 3980
rect 203140 3860 203360 3910
rect 203640 4090 203860 4140
rect 203640 4020 203650 4090
rect 203850 4020 203860 4090
rect 203640 3980 203860 4020
rect 203640 3910 203650 3980
rect 203850 3910 203860 3980
rect 203640 3860 203860 3910
rect 204140 4090 204360 4140
rect 204140 4020 204150 4090
rect 204350 4020 204360 4090
rect 204140 3980 204360 4020
rect 204140 3910 204150 3980
rect 204350 3910 204360 3980
rect 204140 3860 204360 3910
rect 204640 4090 204860 4140
rect 204640 4020 204650 4090
rect 204850 4020 204860 4090
rect 204640 3980 204860 4020
rect 204640 3910 204650 3980
rect 204850 3910 204860 3980
rect 204640 3860 204860 3910
rect 205140 4090 205360 4140
rect 205140 4020 205150 4090
rect 205350 4020 205360 4090
rect 205140 3980 205360 4020
rect 205140 3910 205150 3980
rect 205350 3910 205360 3980
rect 205140 3860 205360 3910
rect 205640 4090 205860 4140
rect 205640 4020 205650 4090
rect 205850 4020 205860 4090
rect 205640 3980 205860 4020
rect 205640 3910 205650 3980
rect 205850 3910 205860 3980
rect 205640 3860 205860 3910
rect 206140 4090 206360 4140
rect 206140 4020 206150 4090
rect 206350 4020 206360 4090
rect 206140 3980 206360 4020
rect 206140 3910 206150 3980
rect 206350 3910 206360 3980
rect 206140 3860 206360 3910
rect 206640 4090 206860 4140
rect 206640 4020 206650 4090
rect 206850 4020 206860 4090
rect 206640 3980 206860 4020
rect 206640 3910 206650 3980
rect 206850 3910 206860 3980
rect 206640 3860 206860 3910
rect 207140 4090 207360 4140
rect 207140 4020 207150 4090
rect 207350 4020 207360 4090
rect 207140 3980 207360 4020
rect 207140 3910 207150 3980
rect 207350 3910 207360 3980
rect 207140 3860 207360 3910
rect 207640 4090 207860 4140
rect 207640 4020 207650 4090
rect 207850 4020 207860 4090
rect 207640 3980 207860 4020
rect 207640 3910 207650 3980
rect 207850 3910 207860 3980
rect 207640 3860 207860 3910
rect 198000 3850 208000 3860
rect 198000 3650 198020 3850
rect 198090 3650 198410 3850
rect 198480 3650 198520 3850
rect 198590 3650 198910 3850
rect 198980 3650 199020 3850
rect 199090 3650 199410 3850
rect 199480 3650 199520 3850
rect 199590 3650 199910 3850
rect 199980 3650 200020 3850
rect 200090 3650 200410 3850
rect 200480 3650 200520 3850
rect 200590 3650 200910 3850
rect 200980 3650 201020 3850
rect 201090 3650 201410 3850
rect 201480 3650 201520 3850
rect 201590 3650 201910 3850
rect 201980 3650 202020 3850
rect 202090 3650 202410 3850
rect 202480 3650 202520 3850
rect 202590 3650 202910 3850
rect 202980 3650 203020 3850
rect 203090 3650 203410 3850
rect 203480 3650 203520 3850
rect 203590 3650 203910 3850
rect 203980 3650 204020 3850
rect 204090 3650 204410 3850
rect 204480 3650 204520 3850
rect 204590 3650 204910 3850
rect 204980 3650 205020 3850
rect 205090 3650 205410 3850
rect 205480 3650 205520 3850
rect 205590 3650 205910 3850
rect 205980 3650 206020 3850
rect 206090 3650 206410 3850
rect 206480 3650 206520 3850
rect 206590 3650 206910 3850
rect 206980 3650 207020 3850
rect 207090 3650 207410 3850
rect 207480 3650 207520 3850
rect 207590 3650 207910 3850
rect 207980 3650 208000 3850
rect 198000 3640 208000 3650
rect 198140 3590 198360 3640
rect 198140 3520 198150 3590
rect 198350 3520 198360 3590
rect 198140 3480 198360 3520
rect 198140 3410 198150 3480
rect 198350 3410 198360 3480
rect 198140 3360 198360 3410
rect 198640 3590 198860 3640
rect 198640 3520 198650 3590
rect 198850 3520 198860 3590
rect 198640 3480 198860 3520
rect 198640 3410 198650 3480
rect 198850 3410 198860 3480
rect 198640 3360 198860 3410
rect 199140 3590 199360 3640
rect 199140 3520 199150 3590
rect 199350 3520 199360 3590
rect 199140 3480 199360 3520
rect 199140 3410 199150 3480
rect 199350 3410 199360 3480
rect 199140 3360 199360 3410
rect 199640 3590 199860 3640
rect 199640 3520 199650 3590
rect 199850 3520 199860 3590
rect 199640 3480 199860 3520
rect 199640 3410 199650 3480
rect 199850 3410 199860 3480
rect 199640 3360 199860 3410
rect 200140 3590 200360 3640
rect 200140 3520 200150 3590
rect 200350 3520 200360 3590
rect 200140 3480 200360 3520
rect 200140 3410 200150 3480
rect 200350 3410 200360 3480
rect 200140 3360 200360 3410
rect 200640 3590 200860 3640
rect 200640 3520 200650 3590
rect 200850 3520 200860 3590
rect 200640 3480 200860 3520
rect 200640 3410 200650 3480
rect 200850 3410 200860 3480
rect 200640 3360 200860 3410
rect 201140 3590 201360 3640
rect 201140 3520 201150 3590
rect 201350 3520 201360 3590
rect 201140 3480 201360 3520
rect 201140 3410 201150 3480
rect 201350 3410 201360 3480
rect 201140 3360 201360 3410
rect 201640 3590 201860 3640
rect 201640 3520 201650 3590
rect 201850 3520 201860 3590
rect 201640 3480 201860 3520
rect 201640 3410 201650 3480
rect 201850 3410 201860 3480
rect 201640 3360 201860 3410
rect 202140 3590 202360 3640
rect 202140 3520 202150 3590
rect 202350 3520 202360 3590
rect 202140 3480 202360 3520
rect 202140 3410 202150 3480
rect 202350 3410 202360 3480
rect 202140 3360 202360 3410
rect 202640 3590 202860 3640
rect 202640 3520 202650 3590
rect 202850 3520 202860 3590
rect 202640 3480 202860 3520
rect 202640 3410 202650 3480
rect 202850 3410 202860 3480
rect 202640 3360 202860 3410
rect 203140 3590 203360 3640
rect 203140 3520 203150 3590
rect 203350 3520 203360 3590
rect 203140 3480 203360 3520
rect 203140 3410 203150 3480
rect 203350 3410 203360 3480
rect 203140 3360 203360 3410
rect 203640 3590 203860 3640
rect 203640 3520 203650 3590
rect 203850 3520 203860 3590
rect 203640 3480 203860 3520
rect 203640 3410 203650 3480
rect 203850 3410 203860 3480
rect 203640 3360 203860 3410
rect 204140 3590 204360 3640
rect 204140 3520 204150 3590
rect 204350 3520 204360 3590
rect 204140 3480 204360 3520
rect 204140 3410 204150 3480
rect 204350 3410 204360 3480
rect 204140 3360 204360 3410
rect 204640 3590 204860 3640
rect 204640 3520 204650 3590
rect 204850 3520 204860 3590
rect 204640 3480 204860 3520
rect 204640 3410 204650 3480
rect 204850 3410 204860 3480
rect 204640 3360 204860 3410
rect 205140 3590 205360 3640
rect 205140 3520 205150 3590
rect 205350 3520 205360 3590
rect 205140 3480 205360 3520
rect 205140 3410 205150 3480
rect 205350 3410 205360 3480
rect 205140 3360 205360 3410
rect 205640 3590 205860 3640
rect 205640 3520 205650 3590
rect 205850 3520 205860 3590
rect 205640 3480 205860 3520
rect 205640 3410 205650 3480
rect 205850 3410 205860 3480
rect 205640 3360 205860 3410
rect 206140 3590 206360 3640
rect 206140 3520 206150 3590
rect 206350 3520 206360 3590
rect 206140 3480 206360 3520
rect 206140 3410 206150 3480
rect 206350 3410 206360 3480
rect 206140 3360 206360 3410
rect 206640 3590 206860 3640
rect 206640 3520 206650 3590
rect 206850 3520 206860 3590
rect 206640 3480 206860 3520
rect 206640 3410 206650 3480
rect 206850 3410 206860 3480
rect 206640 3360 206860 3410
rect 207140 3590 207360 3640
rect 207140 3520 207150 3590
rect 207350 3520 207360 3590
rect 207140 3480 207360 3520
rect 207140 3410 207150 3480
rect 207350 3410 207360 3480
rect 207140 3360 207360 3410
rect 207640 3590 207860 3640
rect 207640 3520 207650 3590
rect 207850 3520 207860 3590
rect 207640 3480 207860 3520
rect 207640 3410 207650 3480
rect 207850 3410 207860 3480
rect 207640 3360 207860 3410
rect 198000 3350 208000 3360
rect 198000 3150 198020 3350
rect 198090 3150 198410 3350
rect 198480 3150 198520 3350
rect 198590 3150 198910 3350
rect 198980 3150 199020 3350
rect 199090 3150 199410 3350
rect 199480 3150 199520 3350
rect 199590 3150 199910 3350
rect 199980 3150 200020 3350
rect 200090 3150 200410 3350
rect 200480 3150 200520 3350
rect 200590 3150 200910 3350
rect 200980 3150 201020 3350
rect 201090 3150 201410 3350
rect 201480 3150 201520 3350
rect 201590 3150 201910 3350
rect 201980 3150 202020 3350
rect 202090 3150 202410 3350
rect 202480 3150 202520 3350
rect 202590 3150 202910 3350
rect 202980 3150 203020 3350
rect 203090 3150 203410 3350
rect 203480 3150 203520 3350
rect 203590 3150 203910 3350
rect 203980 3150 204020 3350
rect 204090 3150 204410 3350
rect 204480 3150 204520 3350
rect 204590 3150 204910 3350
rect 204980 3150 205020 3350
rect 205090 3150 205410 3350
rect 205480 3150 205520 3350
rect 205590 3150 205910 3350
rect 205980 3150 206020 3350
rect 206090 3150 206410 3350
rect 206480 3150 206520 3350
rect 206590 3150 206910 3350
rect 206980 3150 207020 3350
rect 207090 3150 207410 3350
rect 207480 3150 207520 3350
rect 207590 3150 207910 3350
rect 207980 3150 208000 3350
rect 198000 3140 208000 3150
rect 198140 3090 198360 3140
rect 198140 3020 198150 3090
rect 198350 3020 198360 3090
rect 198140 2980 198360 3020
rect 198140 2910 198150 2980
rect 198350 2910 198360 2980
rect 198140 2860 198360 2910
rect 198640 3090 198860 3140
rect 198640 3020 198650 3090
rect 198850 3020 198860 3090
rect 198640 2980 198860 3020
rect 198640 2910 198650 2980
rect 198850 2910 198860 2980
rect 198640 2860 198860 2910
rect 199140 3090 199360 3140
rect 199140 3020 199150 3090
rect 199350 3020 199360 3090
rect 199140 2980 199360 3020
rect 199140 2910 199150 2980
rect 199350 2910 199360 2980
rect 199140 2860 199360 2910
rect 199640 3090 199860 3140
rect 199640 3020 199650 3090
rect 199850 3020 199860 3090
rect 199640 2980 199860 3020
rect 199640 2910 199650 2980
rect 199850 2910 199860 2980
rect 199640 2860 199860 2910
rect 200140 3090 200360 3140
rect 200140 3020 200150 3090
rect 200350 3020 200360 3090
rect 200140 2980 200360 3020
rect 200140 2910 200150 2980
rect 200350 2910 200360 2980
rect 200140 2860 200360 2910
rect 200640 3090 200860 3140
rect 200640 3020 200650 3090
rect 200850 3020 200860 3090
rect 200640 2980 200860 3020
rect 200640 2910 200650 2980
rect 200850 2910 200860 2980
rect 200640 2860 200860 2910
rect 201140 3090 201360 3140
rect 201140 3020 201150 3090
rect 201350 3020 201360 3090
rect 201140 2980 201360 3020
rect 201140 2910 201150 2980
rect 201350 2910 201360 2980
rect 201140 2860 201360 2910
rect 201640 3090 201860 3140
rect 201640 3020 201650 3090
rect 201850 3020 201860 3090
rect 201640 2980 201860 3020
rect 201640 2910 201650 2980
rect 201850 2910 201860 2980
rect 201640 2860 201860 2910
rect 202140 3090 202360 3140
rect 202140 3020 202150 3090
rect 202350 3020 202360 3090
rect 202140 2980 202360 3020
rect 202140 2910 202150 2980
rect 202350 2910 202360 2980
rect 202140 2860 202360 2910
rect 202640 3090 202860 3140
rect 202640 3020 202650 3090
rect 202850 3020 202860 3090
rect 202640 2980 202860 3020
rect 202640 2910 202650 2980
rect 202850 2910 202860 2980
rect 202640 2860 202860 2910
rect 203140 3090 203360 3140
rect 203140 3020 203150 3090
rect 203350 3020 203360 3090
rect 203140 2980 203360 3020
rect 203140 2910 203150 2980
rect 203350 2910 203360 2980
rect 203140 2860 203360 2910
rect 203640 3090 203860 3140
rect 203640 3020 203650 3090
rect 203850 3020 203860 3090
rect 203640 2980 203860 3020
rect 203640 2910 203650 2980
rect 203850 2910 203860 2980
rect 203640 2860 203860 2910
rect 204140 3090 204360 3140
rect 204140 3020 204150 3090
rect 204350 3020 204360 3090
rect 204140 2980 204360 3020
rect 204140 2910 204150 2980
rect 204350 2910 204360 2980
rect 204140 2860 204360 2910
rect 204640 3090 204860 3140
rect 204640 3020 204650 3090
rect 204850 3020 204860 3090
rect 204640 2980 204860 3020
rect 204640 2910 204650 2980
rect 204850 2910 204860 2980
rect 204640 2860 204860 2910
rect 205140 3090 205360 3140
rect 205140 3020 205150 3090
rect 205350 3020 205360 3090
rect 205140 2980 205360 3020
rect 205140 2910 205150 2980
rect 205350 2910 205360 2980
rect 205140 2860 205360 2910
rect 205640 3090 205860 3140
rect 205640 3020 205650 3090
rect 205850 3020 205860 3090
rect 205640 2980 205860 3020
rect 205640 2910 205650 2980
rect 205850 2910 205860 2980
rect 205640 2860 205860 2910
rect 206140 3090 206360 3140
rect 206140 3020 206150 3090
rect 206350 3020 206360 3090
rect 206140 2980 206360 3020
rect 206140 2910 206150 2980
rect 206350 2910 206360 2980
rect 206140 2860 206360 2910
rect 206640 3090 206860 3140
rect 206640 3020 206650 3090
rect 206850 3020 206860 3090
rect 206640 2980 206860 3020
rect 206640 2910 206650 2980
rect 206850 2910 206860 2980
rect 206640 2860 206860 2910
rect 207140 3090 207360 3140
rect 207140 3020 207150 3090
rect 207350 3020 207360 3090
rect 207140 2980 207360 3020
rect 207140 2910 207150 2980
rect 207350 2910 207360 2980
rect 207140 2860 207360 2910
rect 207640 3090 207860 3140
rect 207640 3020 207650 3090
rect 207850 3020 207860 3090
rect 207640 2980 207860 3020
rect 207640 2910 207650 2980
rect 207850 2910 207860 2980
rect 207640 2860 207860 2910
rect 198000 2850 208000 2860
rect 198000 2650 198020 2850
rect 198090 2650 198410 2850
rect 198480 2650 198520 2850
rect 198590 2650 198910 2850
rect 198980 2650 199020 2850
rect 199090 2650 199410 2850
rect 199480 2650 199520 2850
rect 199590 2650 199910 2850
rect 199980 2650 200020 2850
rect 200090 2650 200410 2850
rect 200480 2650 200520 2850
rect 200590 2650 200910 2850
rect 200980 2650 201020 2850
rect 201090 2650 201410 2850
rect 201480 2650 201520 2850
rect 201590 2650 201910 2850
rect 201980 2650 202020 2850
rect 202090 2650 202410 2850
rect 202480 2650 202520 2850
rect 202590 2650 202910 2850
rect 202980 2650 203020 2850
rect 203090 2650 203410 2850
rect 203480 2650 203520 2850
rect 203590 2650 203910 2850
rect 203980 2650 204020 2850
rect 204090 2650 204410 2850
rect 204480 2650 204520 2850
rect 204590 2650 204910 2850
rect 204980 2650 205020 2850
rect 205090 2650 205410 2850
rect 205480 2650 205520 2850
rect 205590 2650 205910 2850
rect 205980 2650 206020 2850
rect 206090 2650 206410 2850
rect 206480 2650 206520 2850
rect 206590 2650 206910 2850
rect 206980 2650 207020 2850
rect 207090 2650 207410 2850
rect 207480 2650 207520 2850
rect 207590 2650 207910 2850
rect 207980 2650 208000 2850
rect 198000 2640 208000 2650
rect 198140 2590 198360 2640
rect 198140 2520 198150 2590
rect 198350 2520 198360 2590
rect 198140 2480 198360 2520
rect 198140 2410 198150 2480
rect 198350 2410 198360 2480
rect 198140 2360 198360 2410
rect 198640 2590 198860 2640
rect 198640 2520 198650 2590
rect 198850 2520 198860 2590
rect 198640 2480 198860 2520
rect 198640 2410 198650 2480
rect 198850 2410 198860 2480
rect 198640 2360 198860 2410
rect 199140 2590 199360 2640
rect 199140 2520 199150 2590
rect 199350 2520 199360 2590
rect 199140 2480 199360 2520
rect 199140 2410 199150 2480
rect 199350 2410 199360 2480
rect 199140 2360 199360 2410
rect 199640 2590 199860 2640
rect 199640 2520 199650 2590
rect 199850 2520 199860 2590
rect 199640 2480 199860 2520
rect 199640 2410 199650 2480
rect 199850 2410 199860 2480
rect 199640 2360 199860 2410
rect 200140 2590 200360 2640
rect 200140 2520 200150 2590
rect 200350 2520 200360 2590
rect 200140 2480 200360 2520
rect 200140 2410 200150 2480
rect 200350 2410 200360 2480
rect 200140 2360 200360 2410
rect 200640 2590 200860 2640
rect 200640 2520 200650 2590
rect 200850 2520 200860 2590
rect 200640 2480 200860 2520
rect 200640 2410 200650 2480
rect 200850 2410 200860 2480
rect 200640 2360 200860 2410
rect 201140 2590 201360 2640
rect 201140 2520 201150 2590
rect 201350 2520 201360 2590
rect 201140 2480 201360 2520
rect 201140 2410 201150 2480
rect 201350 2410 201360 2480
rect 201140 2360 201360 2410
rect 201640 2590 201860 2640
rect 201640 2520 201650 2590
rect 201850 2520 201860 2590
rect 201640 2480 201860 2520
rect 201640 2410 201650 2480
rect 201850 2410 201860 2480
rect 201640 2360 201860 2410
rect 202140 2590 202360 2640
rect 202140 2520 202150 2590
rect 202350 2520 202360 2590
rect 202140 2480 202360 2520
rect 202140 2410 202150 2480
rect 202350 2410 202360 2480
rect 202140 2360 202360 2410
rect 202640 2590 202860 2640
rect 202640 2520 202650 2590
rect 202850 2520 202860 2590
rect 202640 2480 202860 2520
rect 202640 2410 202650 2480
rect 202850 2410 202860 2480
rect 202640 2360 202860 2410
rect 203140 2590 203360 2640
rect 203140 2520 203150 2590
rect 203350 2520 203360 2590
rect 203140 2480 203360 2520
rect 203140 2410 203150 2480
rect 203350 2410 203360 2480
rect 203140 2360 203360 2410
rect 203640 2590 203860 2640
rect 203640 2520 203650 2590
rect 203850 2520 203860 2590
rect 203640 2480 203860 2520
rect 203640 2410 203650 2480
rect 203850 2410 203860 2480
rect 203640 2360 203860 2410
rect 204140 2590 204360 2640
rect 204140 2520 204150 2590
rect 204350 2520 204360 2590
rect 204140 2480 204360 2520
rect 204140 2410 204150 2480
rect 204350 2410 204360 2480
rect 204140 2360 204360 2410
rect 204640 2590 204860 2640
rect 204640 2520 204650 2590
rect 204850 2520 204860 2590
rect 204640 2480 204860 2520
rect 204640 2410 204650 2480
rect 204850 2410 204860 2480
rect 204640 2360 204860 2410
rect 205140 2590 205360 2640
rect 205140 2520 205150 2590
rect 205350 2520 205360 2590
rect 205140 2480 205360 2520
rect 205140 2410 205150 2480
rect 205350 2410 205360 2480
rect 205140 2360 205360 2410
rect 205640 2590 205860 2640
rect 205640 2520 205650 2590
rect 205850 2520 205860 2590
rect 205640 2480 205860 2520
rect 205640 2410 205650 2480
rect 205850 2410 205860 2480
rect 205640 2360 205860 2410
rect 206140 2590 206360 2640
rect 206140 2520 206150 2590
rect 206350 2520 206360 2590
rect 206140 2480 206360 2520
rect 206140 2410 206150 2480
rect 206350 2410 206360 2480
rect 206140 2360 206360 2410
rect 206640 2590 206860 2640
rect 206640 2520 206650 2590
rect 206850 2520 206860 2590
rect 206640 2480 206860 2520
rect 206640 2410 206650 2480
rect 206850 2410 206860 2480
rect 206640 2360 206860 2410
rect 207140 2590 207360 2640
rect 207140 2520 207150 2590
rect 207350 2520 207360 2590
rect 207140 2480 207360 2520
rect 207140 2410 207150 2480
rect 207350 2410 207360 2480
rect 207140 2360 207360 2410
rect 207640 2590 207860 2640
rect 207640 2520 207650 2590
rect 207850 2520 207860 2590
rect 207640 2480 207860 2520
rect 207640 2410 207650 2480
rect 207850 2410 207860 2480
rect 207640 2360 207860 2410
rect 198000 2350 208000 2360
rect 198000 2150 198020 2350
rect 198090 2150 198410 2350
rect 198480 2150 198520 2350
rect 198590 2150 198910 2350
rect 198980 2150 199020 2350
rect 199090 2150 199410 2350
rect 199480 2150 199520 2350
rect 199590 2150 199910 2350
rect 199980 2150 200020 2350
rect 200090 2150 200410 2350
rect 200480 2150 200520 2350
rect 200590 2150 200910 2350
rect 200980 2150 201020 2350
rect 201090 2150 201410 2350
rect 201480 2150 201520 2350
rect 201590 2150 201910 2350
rect 201980 2150 202020 2350
rect 202090 2150 202410 2350
rect 202480 2150 202520 2350
rect 202590 2150 202910 2350
rect 202980 2150 203020 2350
rect 203090 2150 203410 2350
rect 203480 2150 203520 2350
rect 203590 2150 203910 2350
rect 203980 2150 204020 2350
rect 204090 2150 204410 2350
rect 204480 2150 204520 2350
rect 204590 2150 204910 2350
rect 204980 2150 205020 2350
rect 205090 2150 205410 2350
rect 205480 2150 205520 2350
rect 205590 2150 205910 2350
rect 205980 2150 206020 2350
rect 206090 2150 206410 2350
rect 206480 2150 206520 2350
rect 206590 2150 206910 2350
rect 206980 2150 207020 2350
rect 207090 2150 207410 2350
rect 207480 2150 207520 2350
rect 207590 2150 207910 2350
rect 207980 2150 208000 2350
rect 198000 2140 208000 2150
rect 198140 2090 198360 2140
rect 198140 2020 198150 2090
rect 198350 2020 198360 2090
rect 198140 2000 198360 2020
rect 198640 2090 198860 2140
rect 198640 2020 198650 2090
rect 198850 2020 198860 2090
rect 198640 2000 198860 2020
rect 199140 2090 199360 2140
rect 199140 2020 199150 2090
rect 199350 2020 199360 2090
rect 199140 2000 199360 2020
rect 199640 2090 199860 2140
rect 199640 2020 199650 2090
rect 199850 2020 199860 2090
rect 199640 2000 199860 2020
rect 200140 2090 200360 2140
rect 200140 2020 200150 2090
rect 200350 2020 200360 2090
rect 200140 2000 200360 2020
rect 200640 2090 200860 2140
rect 200640 2020 200650 2090
rect 200850 2020 200860 2090
rect 200640 2000 200860 2020
rect 201140 2090 201360 2140
rect 201140 2020 201150 2090
rect 201350 2020 201360 2090
rect 201140 2000 201360 2020
rect 201640 2090 201860 2140
rect 201640 2020 201650 2090
rect 201850 2020 201860 2090
rect 201640 2000 201860 2020
rect 202140 2090 202360 2140
rect 202140 2020 202150 2090
rect 202350 2020 202360 2090
rect 202140 2000 202360 2020
rect 202640 2090 202860 2140
rect 202640 2020 202650 2090
rect 202850 2020 202860 2090
rect 202640 2000 202860 2020
rect 203140 2090 203360 2140
rect 203140 2020 203150 2090
rect 203350 2020 203360 2090
rect 203140 2000 203360 2020
rect 203640 2090 203860 2140
rect 203640 2020 203650 2090
rect 203850 2020 203860 2090
rect 203640 2000 203860 2020
rect 204140 2090 204360 2140
rect 204140 2020 204150 2090
rect 204350 2020 204360 2090
rect 204140 2000 204360 2020
rect 204640 2090 204860 2140
rect 204640 2020 204650 2090
rect 204850 2020 204860 2090
rect 204640 2000 204860 2020
rect 205140 2090 205360 2140
rect 205140 2020 205150 2090
rect 205350 2020 205360 2090
rect 205140 2000 205360 2020
rect 205640 2090 205860 2140
rect 205640 2020 205650 2090
rect 205850 2020 205860 2090
rect 205640 2000 205860 2020
rect 206140 2090 206360 2140
rect 206140 2020 206150 2090
rect 206350 2020 206360 2090
rect 206140 2000 206360 2020
rect 206640 2090 206860 2140
rect 206640 2020 206650 2090
rect 206850 2020 206860 2090
rect 206640 2000 206860 2020
rect 207140 2090 207360 2140
rect 207140 2020 207150 2090
rect 207350 2020 207360 2090
rect 207140 2000 207360 2020
rect 207640 2090 207860 2140
rect 207640 2020 207650 2090
rect 207850 2020 207860 2090
rect 207640 2000 207860 2020
<< via2 >>
rect 250510 135260 250570 135910
rect 171200 119600 172800 121800
rect 222700 119500 224700 121900
rect 128760 86870 128900 87110
rect 129080 86870 129220 87110
rect 128870 86510 129030 86630
rect 129470 67060 129720 67390
<< metal3 >>
rect 250400 135920 250500 136000
rect 250400 135910 250580 135920
rect 250400 135260 250510 135910
rect 250570 135260 250580 135910
rect 250400 135250 250580 135260
rect 250400 135200 250500 135250
rect 16000 121800 22000 124000
rect 68194 123800 73194 124000
rect 68194 122300 73200 123800
rect 68200 122000 73200 122300
rect 16000 116200 16200 121800
rect 21800 116200 22000 121800
rect 16000 116000 22000 116200
rect 120000 121800 126000 124000
rect 165594 122300 170594 124000
rect 170894 122300 173094 124000
rect 173394 122300 175594 124000
rect 175894 122300 180894 124000
rect 217294 122300 222294 124000
rect 222594 122300 224800 124000
rect 225094 122300 227294 124000
rect 227594 122300 232594 124000
rect 318994 122300 323994 124000
rect 324294 122300 326494 124000
rect 326794 122300 328994 124000
rect 329294 122300 334294 124000
rect 413394 122300 418394 124000
rect 465394 123600 470400 124000
rect 465394 122300 465600 123600
rect 120000 116200 120200 121800
rect 125800 116200 126000 121800
rect 120000 116000 126000 116200
rect 166000 121800 170000 122300
rect 166000 115200 166200 121800
rect 169800 115200 170000 121800
rect 171000 121800 173000 122300
rect 171000 119600 171200 121800
rect 172800 119600 173000 121800
rect 171000 119400 173000 119600
rect 166000 115000 170000 115200
rect 173600 119000 175400 122300
rect 218000 121800 222000 122300
rect 173600 114000 181000 119000
rect 218000 115200 218200 121800
rect 221800 115200 222000 121800
rect 222600 121900 224800 122300
rect 222600 119500 222700 121900
rect 224700 119500 224800 121900
rect 222600 119400 224800 119500
rect 218000 115000 222000 115200
rect 225200 114000 227200 122300
rect 465400 121400 465600 122300
rect 469800 121400 470400 123600
rect 510594 123200 515394 124000
rect 510594 122340 515400 123200
rect 520594 122600 525394 124000
rect 520594 122340 525400 122600
rect 465400 121200 470400 121400
rect 510600 122200 515400 122340
rect 510600 116200 510800 122200
rect 515200 116200 515400 122200
rect 510600 115800 515400 116200
rect 520600 122200 525400 122340
rect 566594 122300 571594 124000
rect 520600 116200 520800 122200
rect 525200 116200 525400 122200
rect 520600 115800 525400 116200
rect 0 103000 1700 105242
rect 0 102200 1800 103000
rect 0 100242 1700 102200
rect 582300 97984 584000 102984
rect 130200 87670 132600 87690
rect 130200 87480 130220 87670
rect 128590 87290 130220 87480
rect 132580 87290 132600 87670
rect 128590 87270 132600 87290
rect 133700 87360 136200 87380
rect 128590 87110 128910 87270
rect 133700 87120 133720 87360
rect 128590 86870 128760 87110
rect 128900 86870 128910 87110
rect 128590 86860 128910 86870
rect 129070 87110 133720 87120
rect 129070 86870 129080 87110
rect 129220 86880 133720 87110
rect 136180 86880 136200 87360
rect 129220 86870 136200 86880
rect 129070 86860 136200 86870
rect 128860 86630 129040 86640
rect 128860 86510 128870 86630
rect 129030 86510 129040 86630
rect 128860 86500 129040 86510
rect 128860 86360 129600 86500
rect 0 63842 1660 68642
rect 129460 67400 129600 86360
rect 129460 67390 129730 67400
rect 129460 67060 129470 67390
rect 129720 67060 129730 67390
rect 129460 67050 129730 67060
rect 582340 59784 584000 64584
rect 0 53842 1660 58642
rect 582340 49784 584000 54584
rect 583520 9472 584800 9584
rect 583520 8290 584800 8402
rect 583520 7108 584800 7220
rect 583520 5926 584800 6038
rect 583520 4744 584800 4856
rect 583520 3562 584800 3674
rect 20000 0 20112 400
rect 25400 0 25512 400
rect 30800 0 30912 400
rect 36200 0 36312 400
rect 41600 0 41712 400
rect 47000 0 47112 400
rect 52400 0 52512 400
rect 57800 0 57912 400
rect 63200 0 63312 400
rect 68600 0 68712 400
rect 74000 0 74112 400
rect 79400 0 79512 400
rect 84800 0 84912 400
rect 90200 0 90312 400
rect 95600 0 95712 400
rect 101000 0 101112 400
rect 106400 0 106512 400
rect 111800 0 111912 400
rect 117200 0 117312 400
rect 122600 0 122712 400
rect 128000 0 128112 400
rect 133400 0 133512 400
rect 138800 0 138912 400
rect 144200 0 144312 400
rect 149600 0 149712 400
rect 155000 0 155112 400
rect 160400 0 160512 400
rect 165800 0 165912 400
rect 171200 0 171312 400
rect 176600 0 176712 400
rect 182000 0 182112 400
rect 187400 0 187512 400
rect 192800 0 192912 400
rect 198200 0 198312 400
rect 203600 0 203712 400
rect 209000 0 209112 400
rect 214400 0 214512 400
rect 219800 0 219912 400
rect 225200 0 225312 400
rect 230600 0 230712 400
rect 236000 0 236112 400
rect 241400 0 241512 400
rect 246800 0 246912 400
rect 252200 0 252312 400
rect 257600 0 257712 400
rect 263000 0 263112 400
rect 268400 0 268512 400
rect 273800 0 273912 400
rect 279200 0 279312 400
rect 284600 0 284712 400
rect 290000 0 290112 400
rect 295400 0 295512 400
rect 300800 0 300912 400
rect 306200 0 306312 400
rect 311600 0 311712 400
rect 317000 0 317112 400
rect 322400 0 322512 400
rect 327800 0 327912 400
rect 333200 0 333312 400
rect 338600 0 338712 400
rect 344000 0 344112 400
rect 349400 0 349512 400
rect 354800 0 354912 400
rect 360200 0 360312 400
rect 365600 0 365712 400
rect 371000 0 371112 400
rect 376400 0 376512 400
rect 381800 0 381912 400
rect 387200 0 387312 400
rect 392600 0 392712 400
rect 398000 0 398112 400
rect 403400 0 403512 400
rect 408800 0 408912 400
rect 414200 0 414312 400
rect 419600 0 419712 400
rect 425000 0 425112 400
rect 430400 0 430512 400
rect 435800 0 435912 400
rect 441200 0 441312 400
rect 446600 0 446712 400
rect 452000 0 452112 400
rect 457400 0 457512 400
rect 462800 0 462912 400
rect 468200 0 468312 400
rect 473600 0 473712 400
rect 479000 0 479112 400
rect 484400 0 484512 400
rect 489800 0 489912 400
<< via3 >>
rect 16200 116200 21800 121800
rect 120200 116200 125800 121800
rect 166200 115200 169800 121800
rect 218200 115200 221800 121800
rect 465600 121400 469800 123600
rect 510800 116200 515200 122200
rect 520800 116200 525200 122200
rect 130220 87290 132580 87670
rect 133720 86880 136180 87360
<< metal4 >>
rect 465400 123600 470000 123800
rect 16000 121800 22000 122000
rect 16000 116200 16200 121800
rect 21800 116200 22000 121800
rect 16000 116000 22000 116200
rect 120000 121800 126000 122000
rect 120000 116200 120200 121800
rect 125800 116200 126000 121800
rect 120000 116000 126000 116200
rect 166000 121800 170000 122000
rect 166000 115200 166200 121800
rect 169800 115200 170000 121800
rect 166000 110000 170000 115200
rect 218000 121800 222000 122000
rect 218000 115200 218200 121800
rect 221800 115200 222000 121800
rect 465400 121400 465600 123600
rect 469800 121400 470000 123600
rect 465400 121200 470000 121400
rect 510600 122200 515400 122400
rect 510600 116200 510800 122200
rect 515200 116200 515400 122200
rect 510600 115800 515400 116200
rect 520600 122200 525400 122400
rect 520600 116200 520800 122200
rect 525200 116200 525400 122200
rect 520600 115800 525400 116200
rect 218000 112000 222000 115200
rect 188000 109000 222000 112000
rect 171000 108000 222000 109000
rect 171000 107000 194000 108000
rect 6098 0 13798 800
rect 14458 0 22158 800
rect 24098 0 31798 800
rect 564098 0 571798 800
rect 572458 0 580158 800
<< via4 >>
rect 16200 116200 21800 121800
rect 120200 116200 125800 121800
rect 465600 121400 469800 123600
<< metal5 >>
rect 465400 123600 470000 123800
rect 16000 121800 22000 122000
rect 16000 116200 16200 121800
rect 21800 120000 22000 121800
rect 120000 121800 126000 122000
rect 21800 116200 56000 120000
rect 16000 116000 56000 116200
rect 120000 116200 120200 121800
rect 125800 120000 126000 121800
rect 465400 121400 465600 123600
rect 469800 121400 470000 123600
rect 465400 121200 470000 121400
rect 125800 116200 137000 120000
rect 466000 119800 469400 121200
rect 120000 116000 137000 116200
rect 52000 110000 56000 116000
rect 134000 110000 137000 116000
use RX_top  RX_top_0
timestamp 1662290912
transform 1 0 38000 0 -1 100000
box -37000 -24000 424000 100000
use TX_top  TX_top_0
timestamp 1662290912
transform 1 0 439500 0 -1 83900
box -83500 -40100 132500 83800
use artwork_test_1  artwork_test_1_0
timestamp 1662317594
transform 1 0 253400 0 1 109050
box 0 -99850 99800 -4300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501465
transform 1 0 190000 0 -1 70300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_1
timestamp 1659501465
transform 1 0 192000 0 -1 70300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_2
timestamp 1659501465
transform 1 0 194000 0 -1 70300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_3
timestamp 1659501465
transform 1 0 194000 0 -1 68300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_4
timestamp 1659501465
transform 1 0 194000 0 -1 66300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_154
timestamp 1659501465
transform 1 0 188000 0 -1 70300
box 0 -1700 2000 300
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662263286
transform 1 0 10000 0 -1 122000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_38
timestamp 1662263286
transform 1 0 10000 0 -1 118000
box 0 0 4000 4000
use hash_m1m2m3m4_W20L20_flat  hash_m1m2m3m4_W20L20_flat_93
timestamp 1662263286
transform 1 0 190000 0 -1 70000
box 0 0 4000 4000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660792292
transform 1 0 66000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_1
timestamp 1660792292
transform 1 0 74000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_2
timestamp 1660792292
transform 1 0 82000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_3
timestamp 1660792292
transform 1 0 90000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_4
timestamp 1660792292
transform 1 0 98000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_5
timestamp 1660792292
transform 1 0 106000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_6
timestamp 1660792292
transform 1 0 110000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_7
timestamp 1660792292
transform 1 0 142000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_8
timestamp 1660792292
transform 1 0 150000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_9
timestamp 1660792292
transform 1 0 154000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_10
timestamp 1660792292
transform 1 0 194000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_11
timestamp 1660792292
transform 1 0 186000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_12
timestamp 1660792292
transform 1 0 182000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_13
timestamp 1660792292
transform 1 0 202000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_14
timestamp 1660792292
transform 1 0 206000 0 -1 122000
box 0 0 8000 8000
use hash_m1m2m3m4_W80L80_flat  hash_m1m2m3m4_W80L80_flat_70
timestamp 1660792292
transform 1 0 58000 0 -1 122000
box 0 0 8000 8000
use sky130_fd_pr__nfet_01v8_NLRNVT  sky130_fd_pr__nfet_01v8_NLRNVT_0
timestamp 1662175719
transform 1 0 250611 0 1 135587
box -211 -1187 211 1187
use sky130_fd_pr__res_generic_po_SAMGJE  sky130_fd_pr__res_generic_po_SAMGJE_0
timestamp 1662258694
transform 1 0 128949 0 1 85939
box -469 -939 469 939
<< labels >>
rlabel metal3 s 583520 3562 584800 3674 4 gpio_analog[6]
port 1 nsew
rlabel metal3 s 583520 4744 584800 4856 4 gpio_noesd[6]
port 2 nsew
rlabel metal3 s 582300 97984 584000 102984 4 io_analog[0]
port 3 nsew
rlabel metal3 s 566594 122300 571594 124000 4 io_analog[1]
port 4 nsew
rlabel metal3 s 465394 122300 470394 124000 4 io_analog[2]
port 5 nsew
rlabel metal3 s 413394 122300 418394 124000 4 io_analog[3]
port 6 nsew
rlabel metal3 s 318994 122300 323994 124000 4 io_analog[4]
port 7 nsew
rlabel metal3 s 326794 122300 328994 124000 4 io_clamp_high[0]
port 8 nsew
rlabel metal3 s 324294 122300 326494 124000 4 io_clamp_low[0]
port 9 nsew
rlabel metal3 s 583520 7108 584800 7220 4 io_in[13]
port 10 nsew
rlabel metal3 s 583520 5926 584800 6038 4 io_in_3v3[13]
port 11 nsew
rlabel metal3 s 583520 9472 584800 9584 4 io_oeb[13]
port 12 nsew
rlabel metal3 s 583520 8290 584800 8402 4 io_out[13]
port 13 nsew
rlabel metal3 s 582340 49784 584000 54584 4 vccd1
port 14 nsew
rlabel metal3 s 510594 122340 515394 124000 4 vssa1
port 15 nsew
rlabel metal3 s 173394 122300 175594 124000 4 io_clamp_high[2]
port 16 nsew
rlabel metal3 s 217294 122300 222294 124000 4 io_analog[5]
port 17 nsew
rlabel metal3 s 222594 122300 224794 124000 4 io_clamp_low[1]
port 18 nsew
rlabel metal3 s 170894 122300 173094 124000 4 io_clamp_low[2]
port 19 nsew
rlabel metal3 s 165594 122300 170594 124000 4 io_analog[6]
port 20 nsew
rlabel metal3 s 120194 122300 125194 124000 4 io_analog[7]
port 21 nsew
rlabel metal3 s 68194 122300 73194 124000 4 io_analog[8]
port 22 nsew
rlabel metal3 s 16194 122300 21194 124000 4 io_analog[9]
port 23 nsew
rlabel metal3 s 0 100242 1700 105242 4 io_analog[10]
port 24 nsew
rlabel metal3 s 0 53842 1660 58642 4 vccd2
port 25 nsew
rlabel metal3 s 225094 122300 227294 124000 4 io_clamp_high[1]
port 26 nsew
rlabel metal4 s 572458 0 580158 800 4 vssa1
port 15 nsew
rlabel metal4 s 564098 0 571798 800 4 vdda1
port 120 nsew
rlabel metal4 s 24098 0 31798 800 4 vssa2
port 115 nsew
rlabel metal4 s 14458 0 22158 800 4 vssd2
port 114 nsew
rlabel metal4 s 6098 0 13798 800 4 vdda2
port 113 nsew
rlabel metal3 s 441200 0 441312 400 4 trim[0]
port 112 nsew
rlabel metal3 s 435800 0 435912 400 4 ctln[9]
port 111 nsew
rlabel metal3 s 430400 0 430512 400 4 ctln[8]
port 110 nsew
rlabel metal3 s 425000 0 425112 400 4 ctln[7]
port 109 nsew
rlabel metal3 s 419600 0 419712 400 4 ctln[6]
port 108 nsew
rlabel metal3 s 414200 0 414312 400 4 ctln[5]
port 107 nsew
rlabel metal3 s 408800 0 408912 400 4 ctln[4]
port 106 nsew
rlabel metal3 s 403400 0 403512 400 4 ctln[3]
port 105 nsew
rlabel metal3 s 398000 0 398112 400 4 ctln[2]
port 104 nsew
rlabel metal3 s 392600 0 392712 400 4 ctln[1]
port 103 nsew
rlabel metal3 s 387200 0 387312 400 4 ctln[0]
port 102 nsew
rlabel metal3 s 381800 0 381912 400 4 ctlp[9]
port 101 nsew
rlabel metal3 s 376400 0 376512 400 4 ctlp[8]
port 100 nsew
rlabel metal3 s 371000 0 371112 400 4 ctlp[7]
port 99 nsew
rlabel metal3 s 365600 0 365712 400 4 ctlp[6]
port 98 nsew
rlabel metal3 s 360200 0 360312 400 4 ctlp[5]
port 97 nsew
rlabel metal3 s 354800 0 354912 400 4 ctlp[4]
port 96 nsew
rlabel metal3 s 349400 0 349512 400 4 ctlp[3]
port 95 nsew
rlabel metal3 s 344000 0 344112 400 4 ctlp[2]
port 94 nsew
rlabel metal3 s 338600 0 338712 400 4 ctlp[1]
port 93 nsew
rlabel metal3 s 333200 0 333312 400 4 ctlp[0]
port 92 nsew
rlabel metal3 s 327800 0 327912 400 4 analog_la_in[29]
port 91 nsew
rlabel metal3 s 311600 0 311712 400 4 analog_la_in[28]
port 90 nsew
rlabel metal3 s 306200 0 306312 400 4 analog_la_in[27]
port 89 nsew
rlabel metal3 s 300800 0 300912 400 4 analog_la_in[26]
port 88 nsew
rlabel metal3 s 295400 0 295512 400 4 analog_la_in[25]
port 87 nsew
rlabel metal3 s 489800 0 489912 400 4 trimb[4]
port 86 nsew
rlabel metal3 s 484400 0 484512 400 4 trimb[3]
port 85 nsew
rlabel metal3 s 479000 0 479112 400 4 trimb[2]
port 84 nsew
rlabel metal3 s 473600 0 473712 400 4 trimb[1]
port 83 nsew
rlabel metal3 s 468200 0 468312 400 4 trimb[0]
port 82 nsew
rlabel metal3 s 462800 0 462912 400 4 trim[4]
port 81 nsew
rlabel metal3 s 457400 0 457512 400 4 trim[3]
port 80 nsew
rlabel metal3 s 452000 0 452112 400 4 trim[2]
port 79 nsew
rlabel metal3 s 446600 0 446712 400 4 trim[1]
port 78 nsew
rlabel metal3 s 155000 0 155112 400 4 analog_la_in[19]
port 77 nsew
rlabel metal3 s 149600 0 149712 400 4 analog_la_in[18]
port 76 nsew
rlabel metal3 s 144200 0 144312 400 4 analog_la_in[17]
port 75 nsew
rlabel metal3 s 138800 0 138912 400 4 analog_la_in[16]
port 74 nsew
rlabel metal3 s 133400 0 133512 400 4 analog_la_in[15]
port 73 nsew
rlabel metal3 s 128000 0 128112 400 4 analog_la_in[14]
port 72 nsew
rlabel metal3 s 122600 0 122712 400 4 analog_la_in[13]
port 71 nsew
rlabel metal3 s 117200 0 117312 400 4 analog_la_in[12]
port 70 nsew
rlabel metal3 s 111800 0 111912 400 4 analog_la_in[11]
port 69 nsew
rlabel metal3 s 106400 0 106512 400 4 analog_la_in[10]
port 68 nsew
rlabel metal3 s 101000 0 101112 400 4 analog_la_in[9]
port 67 nsew
rlabel metal3 s 95600 0 95712 400 4 analog_la_in[8]
port 66 nsew
rlabel metal3 s 90200 0 90312 400 4 analog_la_in[7]
port 65 nsew
rlabel metal3 s 84800 0 84912 400 4 analog_la_in[6]
port 64 nsew
rlabel metal3 s 79400 0 79512 400 4 analog_la_in[5]
port 63 nsew
rlabel metal3 s 74000 0 74112 400 4 analog_la_in[4]
port 62 nsew
rlabel metal3 s 68600 0 68712 400 4 analog_la_out[9]
port 61 nsew
rlabel metal3 s 63200 0 63312 400 4 analog_la_out[8]
port 60 nsew
rlabel metal3 s 57800 0 57912 400 4 analog_la_out[7]
port 59 nsew
rlabel metal3 s 52400 0 52512 400 4 analog_la_out[6]
port 58 nsew
rlabel metal3 s 47000 0 47112 400 4 analog_la_out[5]
port 57 nsew
rlabel metal3 s 41600 0 41712 400 4 analog_la_out[4]
port 56 nsew
rlabel metal3 s 36200 0 36312 400 4 analog_la_out[3]
port 55 nsew
rlabel metal3 s 30800 0 30912 400 4 analog_la_out[2]
port 54 nsew
rlabel metal3 s 25400 0 25512 400 4 analog_la_out[1]
port 53 nsew
rlabel metal3 s 20000 0 20112 400 4 analog_la_out[0]
port 52 nsew
rlabel metal3 s 290000 0 290112 400 4 analog_la_in[24]
port 51 nsew
rlabel metal3 s 284600 0 284712 400 4 analog_la_out[29]
port 50 nsew
rlabel metal3 s 279200 0 279312 400 4 analog_la_out[28]
port 49 nsew
rlabel metal3 s 273800 0 273912 400 4 analog_la_out[27]
port 48 nsew
rlabel metal3 s 268400 0 268512 400 4 analog_la_out[26]
port 47 nsew
rlabel metal3 s 263000 0 263112 400 4 analog_la_out[25]
port 46 nsew
rlabel metal3 s 257600 0 257712 400 4 analog_la_out[24]
port 45 nsew
rlabel metal3 s 252200 0 252312 400 4 analog_la_out[23]
port 44 nsew
rlabel metal3 s 246800 0 246912 400 4 analog_la_out[22]
port 43 nsew
rlabel metal3 s 241400 0 241512 400 4 analog_la_out[21]
port 42 nsew
rlabel metal3 s 236000 0 236112 400 4 analog_la_out[20]
port 41 nsew
rlabel metal3 s 230600 0 230712 400 4 analog_la_out[19]
port 40 nsew
rlabel metal3 s 225200 0 225312 400 4 analog_la_out[18]
port 39 nsew
rlabel metal3 s 219800 0 219912 400 4 analog_la_out[17]
port 38 nsew
rlabel metal3 s 214400 0 214512 400 4 analog_la_out[16]
port 37 nsew
rlabel metal3 s 209000 0 209112 400 4 analog_la_out[15]
port 36 nsew
rlabel metal3 s 203600 0 203712 400 4 analog_la_out[14]
port 35 nsew
rlabel metal3 s 198200 0 198312 400 4 analog_la_out[13]
port 34 nsew
rlabel metal3 s 192800 0 192912 400 4 analog_la_out[12]
port 33 nsew
rlabel metal3 s 187400 0 187512 400 4 analog_la_out[11]
port 32 nsew
rlabel metal3 s 182000 0 182112 400 4 analog_la_out[10]
port 31 nsew
rlabel metal3 s 176600 0 176712 400 4 analog_la_in[23]
port 30 nsew
rlabel metal3 s 171200 0 171312 400 4 analog_la_in[22]
port 29 nsew
rlabel metal3 s 165800 0 165912 400 4 analog_la_in[21]
port 28 nsew
rlabel metal3 s 160400 0 160512 400 4 analog_la_in[20]
port 27 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 164000
string path 1929.280 0.000 1929.280 2.000 
<< end >>
