magic
tech sky130B
timestamp 1666835237
<< metal3 >>
rect 1030 1655 1600 1660
rect 1030 1650 2970 1655
rect 1000 1575 2970 1650
rect 1000 1570 1600 1575
rect 1000 1270 1150 1570
rect 1000 1200 2955 1270
rect 1030 1190 2955 1200
rect 1030 1180 1600 1190
rect 1720 570 2800 660
rect 4170 575 4695 655
rect 2190 270 2300 570
rect 4585 270 4695 575
rect 1720 180 2800 270
rect 4170 190 4695 270
rect -580 -40 340 -30
rect -580 -180 120 -40
rect 330 -180 340 -40
rect -580 -190 340 -180
rect -580 -320 340 -310
rect -580 -460 120 -320
rect 330 -460 340 -320
rect -580 -470 340 -460
rect 1720 -790 2800 -700
rect 4170 -770 4695 -690
rect 2190 -1090 2300 -790
rect 4585 -1075 4695 -770
rect 1720 -1180 2800 -1090
rect 4170 -1155 4695 -1075
rect 1490 -1700 2955 -1690
rect 1000 -1770 2955 -1700
rect 1000 -1790 1600 -1770
rect 1000 -2090 1150 -1790
rect 1490 -2090 2955 -2075
rect 1000 -2150 2955 -2090
rect 1030 -2155 2955 -2150
rect 1030 -2180 1600 -2155
<< via3 >>
rect 120 -180 330 -40
rect 120 -460 330 -320
<< metal4 >>
rect 1310 1780 3150 1870
rect 1425 1500 1600 1525
rect 1425 1375 1450 1500
rect 1575 1375 1600 1500
rect 1425 1350 1600 1375
rect 2150 1500 2325 1525
rect 2150 1375 2175 1500
rect 2300 1375 2325 1500
rect 2150 1350 2325 1375
rect 2825 1500 3000 1525
rect 2825 1375 2850 1500
rect 2975 1375 3000 1500
rect 2825 1350 3000 1375
rect -480 910 1190 1040
rect 1315 910 1455 1060
rect 1805 910 1945 1060
rect 3270 910 4940 1040
rect -480 780 1950 910
rect 2510 780 4940 910
rect -480 -1280 -170 780
rect 250 475 425 500
rect 250 350 275 475
rect 400 350 425 475
rect 250 325 425 350
rect 950 475 1125 500
rect 950 350 975 475
rect 1100 350 1125 475
rect 950 325 1125 350
rect 1650 475 1825 500
rect 1650 350 1675 475
rect 1800 350 1825 475
rect 1650 325 1825 350
rect 2650 475 2825 500
rect 2650 350 2675 475
rect 2800 350 2825 475
rect 2650 325 2825 350
rect 3350 475 3525 500
rect 3350 350 3375 475
rect 3500 350 3525 475
rect 3350 325 3525 350
rect 4050 475 4225 500
rect 4050 350 4075 475
rect 4200 350 4225 475
rect 4050 325 4225 350
rect 110 -40 2290 50
rect 2480 30 4350 50
rect 110 -180 120 -40
rect 330 -70 2290 -40
rect 330 -180 1950 -70
rect 110 -190 1950 -180
rect 110 -320 1950 -310
rect 110 -460 120 -320
rect 330 -350 1950 -320
rect 330 -460 1780 -350
rect 110 -530 1780 -460
rect 2080 -430 2290 -70
rect 2590 -150 4350 30
rect 2510 -190 4350 -150
rect 2510 -430 4350 -310
rect 1960 -530 1980 -430
rect 110 -550 1980 -530
rect 2080 -550 4350 -430
rect 250 -875 425 -850
rect 250 -1000 275 -875
rect 400 -1000 425 -875
rect 250 -1025 425 -1000
rect 950 -875 1125 -850
rect 950 -1000 975 -875
rect 1100 -1000 1125 -875
rect 950 -1025 1125 -1000
rect 1625 -875 1800 -850
rect 1625 -1000 1650 -875
rect 1775 -1000 1800 -875
rect 1625 -1025 1800 -1000
rect 2650 -875 2825 -850
rect 2650 -1000 2675 -875
rect 2800 -1000 2825 -875
rect 2650 -1025 2825 -1000
rect 3350 -875 3525 -850
rect 3350 -1000 3375 -875
rect 3500 -1000 3525 -875
rect 3350 -1025 3525 -1000
rect 4025 -875 4200 -850
rect 4025 -1000 4050 -875
rect 4175 -1000 4200 -875
rect 4025 -1025 4200 -1000
rect 4630 -1280 4940 780
rect -480 -1410 1950 -1280
rect 2510 -1410 4940 -1280
rect -480 -1540 1190 -1410
rect 2515 -1560 2655 -1410
rect 3005 -1560 3145 -1410
rect 3270 -1540 4940 -1410
rect 1450 -1875 1625 -1850
rect 1450 -2000 1475 -1875
rect 1600 -2000 1625 -1875
rect 1450 -2025 1625 -2000
rect 2150 -1875 2325 -1850
rect 2150 -2000 2175 -1875
rect 2300 -2000 2325 -1875
rect 2150 -2025 2325 -2000
rect 2850 -1875 3025 -1850
rect 2850 -2000 2875 -1875
rect 3000 -2000 3025 -1875
rect 2850 -2025 3025 -2000
rect 1310 -2370 3150 -2280
<< via4 >>
rect 1450 1375 1575 1500
rect 2175 1375 2300 1500
rect 2850 1375 2975 1500
rect 275 350 400 475
rect 975 350 1100 475
rect 1675 350 1800 475
rect 2675 350 2800 475
rect 3375 350 3500 475
rect 4075 350 4200 475
rect 1780 -530 1960 -350
rect 2410 -150 2590 30
rect 275 -1000 400 -875
rect 975 -1000 1100 -875
rect 1650 -1000 1775 -875
rect 2675 -1000 2800 -875
rect 3375 -1000 3500 -875
rect 4050 -1000 4175 -875
rect 1475 -2000 1600 -1875
rect 2175 -2000 2300 -1875
rect 2875 -2000 3000 -1875
<< metal5 >>
rect -100 1700 1100 1900
rect -100 1400 100 1700
rect 900 1525 1100 1700
rect 3300 1700 4600 1900
rect 3300 1525 3500 1700
rect 900 1500 3500 1525
rect 900 1400 1450 1500
rect -100 1375 1450 1400
rect 1575 1375 2175 1500
rect 2300 1375 2850 1500
rect 2975 1400 3500 1500
rect 4400 1400 4600 1700
rect 2975 1375 4600 1400
rect -100 1350 4600 1375
rect -100 1200 1100 1350
rect -100 500 100 1200
rect 900 500 1100 1200
rect 3300 1200 4600 1350
rect 3300 500 3500 1200
rect 4400 500 4600 1200
rect -100 475 4600 500
rect -100 350 275 475
rect 400 350 975 475
rect 1100 350 1675 475
rect 1800 350 2675 475
rect 2800 350 3375 475
rect 3500 350 4075 475
rect 4200 350 4600 475
rect -100 325 4600 350
rect -100 -850 100 325
rect 900 -850 1100 325
rect 2390 30 2610 50
rect 2390 -130 2410 30
rect 1760 -150 2410 -130
rect 2590 -150 2610 30
rect 1760 -350 2610 -150
rect 1760 -530 1780 -350
rect 1960 -380 2610 -350
rect 1960 -530 1990 -380
rect 1760 -550 1990 -530
rect 3300 -850 3500 325
rect 4400 -850 4600 325
rect -100 -875 4600 -850
rect -100 -1000 275 -875
rect 400 -1000 975 -875
rect 1100 -1000 1650 -875
rect 1775 -1000 2675 -875
rect 2800 -1000 3375 -875
rect 3500 -1000 4050 -875
rect 4175 -1000 4600 -875
rect -100 -1025 4600 -1000
rect -100 -1700 100 -1025
rect 900 -1700 1100 -1025
rect -100 -1850 1100 -1700
rect 3300 -1700 3500 -1025
rect 4400 -1700 4600 -1025
rect 3300 -1850 4600 -1700
rect -100 -1875 4600 -1850
rect -100 -1900 1475 -1875
rect -100 -2200 100 -1900
rect 900 -2000 1475 -1900
rect 1600 -2000 2175 -1875
rect 2300 -2000 2875 -1875
rect 3000 -1900 4600 -1875
rect 3000 -2000 3500 -1900
rect 900 -2025 3500 -2000
rect 900 -2200 1100 -2025
rect -100 -2400 1100 -2200
rect 3300 -2200 3500 -2025
rect 4400 -2200 4600 -1900
rect 3300 -2400 4600 -2200
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_0
timestamp 1659322979
transform 1 0 0 0 1 0
box 0 0 2060 840
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_1
timestamp 1659322979
transform 1 0 2400 0 1 0
box 0 0 2060 840
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_2
timestamp 1659322979
transform 1 0 1200 0 1 1000
box 0 0 2060 840
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_3
timestamp 1659322979
transform 1 0 1200 0 -1 -1500
box 0 0 2060 840
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_4
timestamp 1659322979
transform 1 0 2400 0 -1 -500
box 0 0 2060 840
use RF_nfet_12xW5p0L0p15_fingered_2x  RF_nfet_12xW5p0L0p15_fingered_2x_5
timestamp 1659322979
transform 1 0 0 0 -1 -500
box 0 0 2060 840
<< labels >>
rlabel metal4 1310 1780 3150 1870 1 S1
rlabel metal4 1310 -2370 3150 -2280 1 S2
rlabel metal3 -580 -190 -500 -30 1 IF1
rlabel metal3 -580 -470 -500 -310 1 IF2
rlabel metal3 4590 190 4690 650 1 LO1
rlabel metal3 4590 -1150 4690 -690 1 LO2
rlabel metal3 1000 1200 1100 1650 1 RF1
rlabel metal3 1000 -2150 1100 -1700 1 RF2
rlabel metal5 -100 1700 1100 1900 1 VL
rlabel metal4 -485 780 -170 1040 1 DL
rlabel metal4 4625 -1540 4940 -1280 1 DR
<< end >>
