magic
tech sky130B
magscale 1 2
timestamp 1662605449
<< metal1 >>
rect -1800 -9900 -1300 -9800
rect -1800 -9920 -1680 -9900
rect -1420 -9920 -1300 -9900
rect -1800 -10180 -1700 -9920
rect -1400 -10180 -1300 -9920
rect -1800 -10200 -1680 -10180
rect -1420 -10200 -1300 -10180
rect -1800 -10300 -1300 -10200
<< metal2 >>
rect 30200 9200 33400 9400
rect 30200 7200 30400 9200
rect 33200 7200 33400 9200
rect 34320 7580 34720 7600
rect 34320 7220 34340 7580
rect 34700 7350 34720 7580
rect 34700 7250 35070 7350
rect 34700 7220 34720 7250
rect 34320 7200 34720 7220
rect 30200 7000 33400 7200
rect 30200 1000 30600 7000
rect 31000 1000 31400 7000
rect 31800 1000 32200 7000
rect 32600 1000 33000 7000
rect 34320 6980 34920 7000
rect 34320 6620 34340 6980
rect 34700 6900 34920 6980
rect 34700 6620 34720 6900
rect 34320 6600 34720 6620
rect 34820 6400 34920 6900
rect 34970 6540 35070 7250
rect 34970 6440 35700 6540
rect 34820 6300 35620 6400
rect 34120 6280 34520 6300
rect 34120 5920 34140 6280
rect 34500 6260 34520 6280
rect 34500 6160 35700 6260
rect 34500 5920 34520 6160
rect 34120 5900 34520 5920
rect 34680 6020 35600 6120
rect 34680 5600 34780 6020
rect 34020 5580 34780 5600
rect 34020 5220 34040 5580
rect 34400 5500 34780 5580
rect 34820 5880 35620 5980
rect 34400 5220 34420 5500
rect 34820 5420 34840 5880
rect 35300 5420 35320 5880
rect 34820 5400 35320 5420
rect 34020 5200 34420 5220
rect 30000 800 33200 1000
rect 30000 -1200 30200 800
rect 33000 -1200 33200 800
rect 30000 -1400 33200 -1200
<< via2 >>
rect 30400 7200 33200 9200
rect 34340 7220 34700 7580
rect 34340 6620 34700 6980
rect 34140 5920 34500 6280
rect 34040 5220 34400 5580
rect 34840 5420 35300 5880
rect 30200 -1200 33000 800
<< metal3 >>
rect 30200 9200 33400 9400
rect 17120 6900 21400 7700
rect 30200 7200 30400 9200
rect 33200 7200 33400 9200
rect 34420 8980 35220 9400
rect 30200 7000 33400 7200
rect 33940 8960 35220 8980
rect 33940 8400 34440 8960
rect 35200 8400 35220 8960
rect 33940 8380 35220 8400
rect 17120 6700 18200 6900
rect 33940 6300 34240 8380
rect 34320 7580 34720 7600
rect 34320 7220 34340 7580
rect 34700 7220 34720 7580
rect 34320 7200 34720 7220
rect 34320 6980 34720 7000
rect 34320 6620 34340 6980
rect 34700 6620 34720 6980
rect 34320 6600 34720 6620
rect 33940 6280 34520 6300
rect 33940 5920 34140 6280
rect 34500 5920 34520 6280
rect 33940 5900 34520 5920
rect 34820 5880 35320 5900
rect 28600 5000 31800 5800
rect 34020 5580 34420 5600
rect 34020 5220 34040 5580
rect 34400 5220 34420 5580
rect 34820 5420 34840 5880
rect 35300 5420 35320 5880
rect 34820 5400 35320 5420
rect 34020 5200 34420 5220
rect 29600 4500 30200 4600
rect 26540 4480 30200 4500
rect 26540 4140 26560 4480
rect 28040 4140 30200 4480
rect 26540 4120 30200 4140
rect 26540 3860 30400 3880
rect 26540 3520 26560 3860
rect 28040 3520 30400 3860
rect 26540 3500 30400 3520
rect 29800 3400 30400 3500
rect 31000 3400 31800 5000
rect 28600 2200 30200 3000
rect 31000 2600 34600 3400
rect 29600 1400 34600 2200
rect 14200 1200 18200 1300
rect 14200 -1000 14300 1200
rect 16900 1100 18200 1200
rect 16900 300 21600 1100
rect 30020 800 33220 1000
rect 16900 -1000 17000 300
rect 14200 -1100 17000 -1000
rect 30020 -1200 30200 800
rect 33020 700 33220 800
rect 33020 -300 38720 700
rect 33020 -1200 33220 -300
rect 30020 -1400 33220 -1200
rect 36720 -1300 38720 -300
<< via3 >>
rect 30400 7200 33200 9200
rect 34440 8400 35200 8960
rect 34340 7220 34700 7580
rect 34340 6620 34700 6980
rect 34040 5220 34400 5580
rect 34840 5420 35300 5880
rect 26560 4140 28040 4480
rect 26560 3520 28040 3860
rect 14300 -1000 16900 1200
rect 30220 -1200 33000 800
rect 33000 -1200 33020 800
<< metal4 >>
rect 6720 22700 20720 24700
rect 17720 11700 20720 22700
rect 30620 17600 32720 17700
rect 30620 14800 30720 17600
rect 32620 14800 32720 17600
rect 30620 12200 32720 14800
rect 17720 10500 29720 11700
rect 17720 9700 29800 10500
rect 30620 10100 34020 12200
rect 22200 8240 25400 9500
rect 21980 8100 25660 8240
rect 28600 5900 29800 9700
rect 30200 9200 33400 9400
rect 30200 7200 30400 9200
rect 33200 7200 33400 9200
rect 33520 7600 34020 10100
rect 34420 8960 35220 9400
rect 34420 8400 34440 8960
rect 35200 8400 35220 8960
rect 34420 8380 35220 8400
rect 33520 7580 34720 7600
rect 33520 7220 34340 7580
rect 34700 7220 34720 7580
rect 33520 7200 34720 7220
rect 30200 7000 33400 7200
rect 33520 6980 34720 7000
rect 33520 6620 34340 6980
rect 34700 6620 34720 6980
rect 33520 6600 34720 6620
rect 33520 6200 33920 6600
rect 32400 5800 33920 6200
rect 34820 5880 35320 5900
rect 32400 4800 32800 5800
rect 29800 4600 32800 4800
rect 29600 4400 32800 4600
rect 33000 5580 34420 5600
rect 33000 5220 34040 5580
rect 34400 5220 34420 5580
rect 33000 5200 34420 5220
rect 34820 5420 34840 5880
rect 35300 5420 35320 5880
rect 34820 5200 35320 5420
rect 29600 4200 30200 4400
rect 33000 4200 33400 5200
rect 30400 3800 33400 4200
rect 29800 3400 30800 3800
rect 17800 1900 18400 3300
rect 11400 1200 17000 1300
rect 11400 -1000 14300 1200
rect 16900 -1000 17000 1200
rect 11400 -1100 17000 -1000
rect 17800 -2100 19000 1900
rect 30000 800 33220 1000
rect 22200 -1500 25400 -100
rect 30000 -1200 30200 800
rect 33020 -1200 33220 800
rect 30000 -1400 33220 -1200
rect 34800 -1300 35400 5200
rect 34220 -1400 36220 -1300
rect 17800 -10700 19400 -2100
rect 34220 -3200 34320 -1400
rect 36120 -3200 36220 -1400
rect 34220 -3300 36220 -3200
rect 25820 -10700 27920 -10681
rect 17720 -10793 27920 -10700
rect 17720 -12569 26032 -10793
rect 27808 -12569 27920 -10793
rect 17720 -12700 27920 -12569
<< via4 >>
rect 30720 14800 32620 17600
rect 30400 7200 33200 9200
rect 30200 -1200 30220 800
rect 30220 -1200 33020 800
rect 34320 -3200 36120 -1400
rect 26032 -12569 27808 -10793
<< metal5 >>
rect 31720 20500 32620 21100
rect 29720 18700 32620 20500
rect 28020 17700 32620 18700
rect 28020 17600 32720 17700
rect 28020 17000 30720 17600
rect 26320 15700 30720 17000
rect 24720 14800 30720 15700
rect 32620 14800 32720 17600
rect 24720 14700 32720 14800
rect 20200 8700 28200 9500
rect 20200 8300 20600 8700
rect 21000 8300 21400 8700
rect 22200 8500 25400 8700
rect 26200 8300 26600 8700
rect 27000 8300 27400 8700
rect 27800 8300 28200 8700
rect 30000 9200 33400 9400
rect 30000 8300 30400 9200
rect 28400 7200 30400 8300
rect 33200 7200 33400 9200
rect 28400 6900 33400 7200
rect 28400 800 33220 1100
rect 20200 -700 20600 -100
rect 21000 -700 21400 -100
rect 22200 -700 25400 -500
rect 26200 -700 26600 -100
rect 27000 -700 27400 -100
rect 27800 -200 28200 -100
rect 28400 -200 30200 800
rect 27800 -700 30200 -200
rect 20200 -1200 30200 -700
rect 33020 -1200 33220 800
rect 20200 -1400 33220 -1200
rect 34220 -1400 36220 -1300
rect 20200 -1500 28200 -1400
rect 34220 -3200 34320 -1400
rect 36120 -3200 36220 -1400
rect 34220 -3300 36220 -3200
tri 24168 -5300 26168 -3300 se
rect 26168 -5300 47272 -3300
tri 47272 -5300 49272 -3300 sw
tri 21568 -7900 24168 -5300 se
rect 24168 -5900 26396 -5300
tri 26396 -5900 26996 -5300 nw
tri 46444 -5900 47044 -5300 ne
rect 47044 -5900 49272 -5300
rect 24168 -6749 25547 -5900
tri 25547 -6749 26396 -5900 nw
tri 26396 -6749 27245 -5900 se
rect 27245 -6749 46195 -5900
tri 46195 -6749 47044 -5900 sw
tri 47044 -6749 47893 -5900 ne
rect 47893 -6749 49272 -5900
rect 24168 -7051 25245 -6749
tri 25245 -7051 25547 -6749 nw
tri 26094 -7051 26396 -6749 se
rect 26396 -6976 47044 -6749
tri 47044 -6976 47271 -6749 sw
tri 47893 -6976 48120 -6749 ne
rect 48120 -6976 49272 -6749
tri 49272 -6976 50948 -5300 sw
rect 26396 -7051 47271 -6976
rect 24168 -7900 24396 -7051
tri 24396 -7900 25245 -7051 nw
tri 25245 -7900 26094 -7051 se
rect 26094 -7825 47271 -7051
tri 47271 -7825 48120 -6976 sw
tri 48120 -7825 48969 -6976 ne
rect 48969 -7825 50948 -6976
rect 26094 -7900 48120 -7825
tri 20720 -8748 21568 -7900 se
rect 21568 -8748 23547 -7900
rect 20720 -8749 23547 -8748
tri 23547 -8749 24396 -7900 nw
tri 24396 -8749 25245 -7900 se
rect 25245 -8500 27473 -7900
tri 27473 -8500 28073 -7900 nw
tri 45367 -8500 45967 -7900 ne
rect 45967 -8053 48120 -7900
tri 48120 -8053 48348 -7825 sw
tri 48969 -8053 49197 -7825 ne
rect 49197 -8053 50948 -7825
rect 45967 -8500 48348 -8053
rect 25245 -8749 26624 -8500
rect 20720 -14385 22720 -8749
tri 22720 -9576 23547 -8749 nw
tri 23569 -9576 24396 -8749 se
rect 24396 -9349 26624 -8749
tri 26624 -9349 27473 -8500 nw
tri 27473 -9349 28322 -8500 se
rect 28322 -8902 45118 -8500
tri 45118 -8902 45520 -8500 sw
tri 45967 -8902 46369 -8500 ne
rect 46369 -8902 48348 -8500
tri 48348 -8902 49197 -8053 sw
tri 49197 -8902 50046 -8053 ne
rect 50046 -8748 50948 -8053
tri 50948 -8748 52720 -6976 sw
rect 50046 -8902 52720 -8748
rect 28322 -9349 45520 -8902
rect 24396 -9576 26322 -9349
tri 23320 -9825 23569 -9576 se
rect 23569 -9651 26322 -9576
tri 26322 -9651 26624 -9349 nw
tri 27171 -9651 27473 -9349 se
rect 27473 -9651 45520 -9349
rect 23569 -9825 25473 -9651
rect 23320 -10500 25473 -9825
tri 25473 -10500 26322 -9651 nw
tri 26322 -10500 27171 -9651 se
rect 27171 -9751 45520 -9651
tri 45520 -9751 46369 -8902 sw
tri 46369 -9751 47218 -8902 ne
rect 47218 -9576 49197 -8902
tri 49197 -9576 49871 -8902 sw
tri 50046 -9576 50720 -8902 ne
rect 47218 -9751 49871 -9576
rect 27171 -10500 46369 -9751
tri 46369 -10500 47118 -9751 sw
tri 47218 -10500 47967 -9751 ne
rect 47967 -9825 49871 -9751
tri 49871 -9825 50120 -9576 sw
rect 50720 -9700 52720 -8902
rect 47967 -10500 50120 -9825
rect 23320 -13537 25320 -10500
tri 25320 -10653 25473 -10500 nw
tri 26141 -10681 26322 -10500 se
rect 26322 -10681 27920 -10500
rect 25920 -10793 27920 -10681
rect 25920 -12569 26032 -10793
rect 27808 -12569 27920 -10793
tri 27920 -11730 29150 -10500 nw
tri 44290 -11730 45520 -10500 ne
rect 45520 -10902 47118 -10500
tri 47118 -10902 47520 -10500 sw
tri 47967 -10653 48120 -10500 ne
rect 25920 -12681 27920 -12569
tri 22720 -14385 23320 -13785 sw
tri 23320 -14385 24168 -13537 ne
rect 24168 -14385 25320 -13537
rect 20720 -14614 23320 -14385
tri 20720 -16614 22720 -14614 ne
rect 22720 -14700 23320 -14614
tri 23320 -14700 23635 -14385 sw
tri 24168 -14700 24483 -14385 ne
rect 24483 -14700 25320 -14385
tri 25320 -14700 27312 -12708 sw
tri 43528 -14700 45520 -12708 se
rect 45520 -13537 47520 -10902
rect 45520 -14385 46672 -13537
tri 46672 -14385 47520 -13537 nw
tri 47520 -14385 48120 -13785 se
rect 48120 -14385 50120 -10500
rect 45520 -14700 46357 -14385
tri 46357 -14700 46672 -14385 nw
tri 47205 -14700 47520 -14385 se
rect 47520 -14614 50120 -14385
rect 47520 -14700 50034 -14614
tri 50034 -14700 50120 -14614 nw
rect 22720 -15537 23635 -14700
tri 23635 -15537 24472 -14700 sw
tri 24483 -15537 25320 -14700 ne
rect 25320 -15537 45509 -14700
rect 22720 -16385 24472 -15537
tri 24472 -16385 25320 -15537 sw
tri 25320 -16385 26168 -15537 ne
rect 26168 -15548 45509 -15537
tri 45509 -15548 46357 -14700 nw
tri 46357 -15548 47205 -14700 se
rect 47205 -15548 47434 -14700
rect 26168 -15852 45205 -15548
tri 45205 -15852 45509 -15548 nw
tri 46053 -15852 46357 -15548 se
rect 46357 -15852 47434 -15548
rect 26168 -16385 44357 -15852
rect 22720 -16614 25320 -16385
tri 22720 -19214 25320 -16614 ne
tri 25320 -16700 25635 -16385 sw
tri 26168 -16700 26483 -16385 ne
rect 26483 -16700 44357 -16385
tri 44357 -16700 45205 -15852 nw
tri 45205 -16700 46053 -15852 se
rect 46053 -16700 47434 -15852
rect 25320 -17300 25635 -16700
tri 25635 -17300 26235 -16700 sw
tri 44605 -17300 45205 -16700 se
rect 45205 -17300 47434 -16700
tri 47434 -17300 50034 -14700 nw
rect 25320 -19214 45434 -17300
tri 25320 -19300 25406 -19214 ne
rect 25406 -19300 45434 -19214
tri 45434 -19300 47434 -17300 nw
use MIXER_5G_core  MIXER_5G_core_0
timestamp 1662605449
transform 1 0 19360 0 1 4500
box -1160 -4800 9880 3800
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1659501465
transform 0 1 54420 1 0 -15300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_1
timestamp 1659501465
transform 0 1 50420 1 0 -21300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_4
timestamp 1659501465
transform 0 1 52420 1 0 -3300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_10
timestamp 1659501465
transform 0 1 52420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_11
timestamp 1659501465
transform 0 1 50420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_12
timestamp 1659501465
transform 0 1 48420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_13
timestamp 1659501465
transform 0 1 46420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_14
timestamp 1659501465
transform 0 1 44420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_15
timestamp 1659501465
transform 0 1 42420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_16
timestamp 1659501465
transform 0 1 40420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_17
timestamp 1659501465
transform 0 1 38420 1 0 -1300
box 0 -1700 2000 300
use hash_m1m2m3m4_W10L10_flat  hash_m1m2m3m4_W10L10_flat_18
timestamp 1659501465
transform 0 1 54420 1 0 -17300
box 0 -1700 2000 300
use mixer_biasgen  mixer_biasgen_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1662239336
transform 1 0 36020 0 -1 6080
box -420 -2040 9600 1680
use octa_ind_700p_thinner  octa_ind_700p_thinner_1 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1662238829
transform -1 0 14420 0 -1 22700
box -17300 -8000 14700 8000
<< end >>
