magic
tech sky130B
magscale 1 2
timestamp 1660522229
<< error_p >>
rect -47842 -11958 -47800 -11680
rect -48120 -12000 -47800 -11958
rect -47616 -12226 -47574 -12184
<< metal4 >>
rect -48400 -24112 -34600 -24000
rect -48400 -27888 -48288 -24112
rect -44512 -27888 -38488 -24112
rect -34712 -27888 -34600 -24112
rect -48400 -28000 -34600 -27888
<< via4 >>
rect -48288 -27888 -44512 -24112
rect -38488 -27888 -34712 -24112
<< metal5 >>
rect -32800 400 -11620 3000
rect -35200 -1000 -11620 400
tri -11620 -1000 -7620 3000 sw
rect -35200 -1600 -31923 -1000
tri -31923 -1600 -31323 -1000 nw
tri -13277 -1600 -12677 -1000 ne
rect -12677 -1600 -7620 -1000
rect -35200 -2449 -32772 -1600
tri -32772 -2449 -31923 -1600 nw
tri -31923 -2449 -31074 -1600 se
rect -31074 -2449 -13526 -1600
tri -13526 -2449 -12677 -1600 sw
tri -12677 -2449 -11828 -1600 ne
rect -11828 -2449 -7620 -1600
rect -35200 -2800 -33621 -2449
rect -36800 -3298 -33621 -2800
tri -33621 -3298 -32772 -2449 nw
tri -32772 -3298 -31923 -2449 se
rect -31923 -3298 -12677 -2449
tri -12677 -3298 -11828 -2449 sw
tri -11828 -3298 -10979 -2449 ne
rect -10979 -3298 -7620 -2449
rect -36800 -3902 -34225 -3298
tri -34225 -3902 -33621 -3298 nw
tri -33376 -3902 -32772 -3298 se
rect -32772 -3902 -11828 -3298
tri -11828 -3902 -11224 -3298 sw
tri -10979 -3902 -10375 -3298 ne
rect -10375 -3902 -7620 -3298
rect -36800 -4751 -35074 -3902
tri -35074 -4751 -34225 -3902 nw
tri -34225 -4751 -33376 -3902 se
rect -33376 -4751 -11224 -3902
tri -11224 -4751 -10375 -3902 sw
tri -10375 -4751 -9526 -3902 ne
rect -9526 -4751 -7620 -3902
rect -36800 -5400 -35923 -4751
rect -39600 -5600 -35923 -5400
tri -35923 -5600 -35074 -4751 nw
tri -35074 -5600 -34225 -4751 se
rect -34225 -5600 -10375 -4751
tri -10375 -5600 -9526 -4751 sw
tri -9526 -5600 -8677 -4751 ne
rect -8677 -5600 -7620 -4751
tri -7620 -5600 -3020 -1000 sw
rect -39600 -6449 -36772 -5600
tri -36772 -6449 -35923 -5600 nw
tri -35923 -6449 -35074 -5600 se
rect -39600 -7298 -37621 -6449
tri -37621 -7298 -36772 -6449 nw
tri -36772 -7298 -35923 -6449 se
rect -35923 -7298 -35074 -6449
rect -39600 -8028 -38351 -7298
tri -38351 -8028 -37621 -7298 nw
tri -37502 -8028 -36772 -7298 se
rect -36772 -8028 -35074 -7298
rect -39600 -8400 -39200 -8028
rect -43600 -8877 -39200 -8400
tri -39200 -8877 -38351 -8028 nw
tri -38351 -8877 -37502 -8028 se
rect -37502 -8877 -35074 -8028
rect -43600 -9726 -40049 -8877
tri -40049 -9726 -39200 -8877 nw
tri -39200 -9726 -38351 -8877 se
rect -38351 -9726 -35074 -8877
rect -43600 -10575 -40898 -9726
tri -40898 -10575 -40049 -9726 nw
tri -40049 -10575 -39200 -9726 se
rect -39200 -10575 -35074 -9726
rect -43600 -11000 -41580 -10575
rect -57600 -11257 -41580 -11000
tri -41580 -11257 -40898 -10575 nw
tri -40731 -11257 -40049 -10575 se
rect -40049 -11257 -35074 -10575
tri -35074 -11257 -29417 -5600 nw
tri -15183 -11257 -9526 -5600 ne
tri -9526 -6449 -8677 -5600 sw
tri -8677 -6449 -7828 -5600 ne
rect -7828 -6449 -3020 -5600
rect -9526 -7298 -8677 -6449
tri -8677 -7298 -7828 -6449 sw
tri -7828 -7298 -6979 -6449 ne
rect -6979 -7298 -3020 -6449
rect -9526 -8028 -7828 -7298
tri -7828 -8028 -7098 -7298 sw
tri -6979 -8028 -6249 -7298 ne
rect -6249 -8028 -3020 -7298
rect -9526 -8877 -7098 -8028
tri -7098 -8877 -6249 -8028 sw
tri -6249 -8877 -5400 -8028 ne
rect -5400 -8877 -3020 -8028
rect -9526 -9726 -6249 -8877
tri -6249 -9726 -5400 -8877 sw
tri -5400 -9726 -4551 -8877 ne
rect -4551 -9726 -3020 -8877
tri -3020 -9726 1106 -5600 sw
rect -9526 -10575 -5400 -9726
tri -5400 -10575 -4551 -9726 sw
tri -4551 -10575 -3702 -9726 ne
rect -3702 -10575 1106 -9726
rect -9526 -11257 -4551 -10575
rect -57600 -11958 -42323 -11257
rect -57600 -12000 -47842 -11958
tri -47842 -12000 -47800 -11958 nw
rect -47800 -12000 -42323 -11958
tri -42323 -12000 -41580 -11257 nw
tri -41474 -12000 -40731 -11257 se
rect -40731 -12000 -39200 -11257
rect -57600 -12849 -43172 -12000
tri -43172 -12849 -42323 -12000 nw
tri -42323 -12849 -41474 -12000 se
rect -41474 -12849 -39200 -12000
rect -57600 -16000 -43800 -12849
tri -43800 -13477 -43172 -12849 nw
tri -42951 -13477 -42323 -12849 se
rect -42323 -13477 -39200 -12849
tri -43200 -13726 -42951 -13477 se
rect -42951 -13726 -39200 -13477
rect -57600 -24112 -44400 -24000
rect -57600 -27888 -48288 -24112
rect -44512 -27888 -44400 -24112
rect -57600 -28000 -44400 -27888
rect -43200 -28470 -39200 -13726
tri -39200 -15383 -35074 -11257 nw
tri -9526 -15383 -5400 -11257 ne
rect -5400 -11424 -4551 -11257
tri -4551 -11424 -3702 -10575 sw
tri -3702 -11424 -2853 -10575 ne
rect -2853 -11424 1106 -10575
rect -5400 -12028 -3702 -11424
tri -3702 -12028 -3098 -11424 sw
tri -2853 -12028 -2249 -11424 ne
rect -2249 -11820 1106 -11424
tri 1106 -11820 3200 -9726 sw
rect -2249 -12028 3200 -11820
rect -5400 -12877 -3098 -12028
tri -3098 -12877 -2249 -12028 sw
tri -2249 -12877 -1400 -12028 ne
rect -1400 -12877 3200 -12028
rect -5400 -13726 -2249 -12877
tri -2249 -13726 -1400 -12877 sw
tri -1400 -13477 -800 -12877 ne
rect -38600 -24112 -34600 -24000
tri -39200 -28470 -38600 -27870 sw
rect -38600 -27888 -38488 -24112
rect -34712 -27888 -34600 -24112
rect -38600 -28000 -34600 -27888
tri -38222 -28470 -37752 -28000 ne
rect -37752 -28470 -34600 -28000
rect -43200 -29318 -38600 -28470
tri -38600 -29318 -37752 -28470 sw
tri -37752 -29318 -36904 -28470 ne
rect -36904 -29318 -34600 -28470
rect -43200 -29527 -37752 -29318
tri -43200 -34400 -38327 -29527 ne
rect -38327 -29926 -37752 -29527
tri -37752 -29926 -37144 -29318 sw
tri -36904 -29926 -36296 -29318 ne
rect -36296 -29926 -34600 -29318
rect -38327 -30774 -37144 -29926
tri -37144 -30774 -36296 -29926 sw
tri -36296 -30774 -35448 -29926 ne
rect -35448 -30774 -34600 -29926
rect -38327 -31622 -36296 -30774
tri -36296 -31622 -35448 -30774 sw
tri -35448 -31622 -34600 -30774 ne
tri -34600 -31622 -28943 -25965 sw
tri -7435 -28000 -5400 -25965 se
rect -5400 -27622 -1400 -13726
rect -5400 -28000 -2248 -27622
tri -8178 -28743 -7435 -28000 se
rect -7435 -28470 -2248 -28000
tri -2248 -28470 -1400 -27622 nw
tri -1400 -28470 -800 -27870 se
rect -800 -28470 3200 -12877
rect -7435 -28743 -2521 -28470
tri -2521 -28743 -2248 -28470 nw
tri -1673 -28743 -1400 -28470 se
rect -1400 -28743 3200 -28470
tri -11057 -31622 -8178 -28743 se
rect -8178 -29591 -3369 -28743
tri -3369 -29591 -2521 -28743 nw
tri -2521 -29591 -1673 -28743 se
rect -1673 -29527 3200 -28743
rect -1673 -29591 -800 -29527
rect -8178 -29926 -3704 -29591
tri -3704 -29926 -3369 -29591 nw
tri -2856 -29926 -2521 -29591 se
rect -2521 -29926 -800 -29591
rect -8178 -30774 -4552 -29926
tri -4552 -30774 -3704 -29926 nw
tri -3704 -30774 -2856 -29926 se
rect -2856 -30774 -800 -29926
rect -8178 -31622 -5400 -30774
tri -5400 -31622 -4552 -30774 nw
tri -4552 -31622 -3704 -30774 se
rect -3704 -31622 -800 -30774
rect -38327 -32470 -35448 -31622
tri -35448 -32470 -34600 -31622 sw
tri -34600 -32470 -33752 -31622 ne
rect -33752 -32470 -28943 -31622
rect -38327 -33318 -34600 -32470
tri -34600 -33318 -33752 -32470 sw
tri -33752 -33318 -32904 -32470 ne
rect -32904 -33318 -28943 -32470
rect -38327 -33552 -33752 -33318
tri -33752 -33552 -33518 -33318 sw
tri -32904 -33552 -32670 -33318 ne
rect -32670 -33552 -28943 -33318
rect -38327 -34400 -33518 -33552
tri -33518 -34400 -32670 -33552 sw
tri -32670 -34400 -31822 -33552 ne
rect -31822 -34400 -28943 -33552
tri -28943 -34400 -26165 -31622 sw
tri -13835 -34400 -11057 -31622 se
rect -11057 -32470 -6248 -31622
tri -6248 -32470 -5400 -31622 nw
tri -5400 -32470 -4552 -31622 se
rect -4552 -32470 -800 -31622
rect -11057 -33318 -7096 -32470
tri -7096 -33318 -6248 -32470 nw
tri -6248 -33318 -5400 -32470 se
rect -5400 -33318 -800 -32470
rect -11057 -33552 -7330 -33318
tri -7330 -33552 -7096 -33318 nw
tri -6482 -33552 -6248 -33318 se
rect -6248 -33527 -800 -33318
tri -800 -33527 3200 -29527 nw
rect -6248 -33552 -5400 -33527
rect -11057 -34400 -8178 -33552
tri -8178 -34400 -7330 -33552 nw
tri -7330 -34400 -6482 -33552 se
rect -6482 -34400 -5400 -33552
tri -38327 -39000 -33727 -34400 ne
rect -33727 -35248 -32670 -34400
tri -32670 -35248 -31822 -34400 sw
tri -31822 -35248 -30974 -34400 ne
rect -30974 -35248 -9026 -34400
tri -9026 -35248 -8178 -34400 nw
tri -8178 -35248 -7330 -34400 se
rect -7330 -35248 -5400 -34400
rect -33727 -36096 -31822 -35248
tri -31822 -36096 -30974 -35248 sw
tri -30974 -36096 -30126 -35248 ne
rect -30126 -36096 -9874 -35248
tri -9874 -36096 -9026 -35248 nw
tri -9026 -36096 -8178 -35248 se
rect -8178 -36096 -5400 -35248
rect -33727 -36704 -30974 -36096
tri -30974 -36704 -30366 -36096 sw
tri -30126 -36704 -29518 -36096 ne
rect -29518 -36704 -10482 -36096
tri -10482 -36704 -9874 -36096 nw
tri -9634 -36704 -9026 -36096 se
rect -9026 -36704 -5400 -36096
rect -33727 -37552 -30366 -36704
tri -30366 -37552 -29518 -36704 sw
tri -29518 -37552 -28670 -36704 ne
rect -28670 -37552 -11330 -36704
tri -11330 -37552 -10482 -36704 nw
tri -10482 -37552 -9634 -36704 se
rect -9634 -37552 -5400 -36704
rect -33727 -38400 -29518 -37552
tri -29518 -38400 -28670 -37552 sw
tri -28670 -38400 -27822 -37552 ne
rect -27822 -38400 -12178 -37552
tri -12178 -38400 -11330 -37552 nw
tri -11330 -38400 -10482 -37552 se
rect -10482 -38127 -5400 -37552
tri -5400 -38127 -800 -33527 nw
rect -10482 -38400 -10273 -38127
rect -33727 -39000 -28670 -38400
tri -28670 -39000 -28070 -38400 sw
tri -11930 -39000 -11330 -38400 se
rect -11330 -39000 -10273 -38400
tri -33727 -43000 -29727 -39000 ne
rect -29727 -43000 -10273 -39000
tri -10273 -43000 -5400 -38127 nw
<< end >>
