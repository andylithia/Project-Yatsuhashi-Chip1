magic
tech sky130B
magscale 1 2
timestamp 1660736647
<< metal2 >>
rect -508 2208 -381 2680
rect -2020 2100 -1760 2140
rect -2020 2020 -1980 2100
rect -1860 2020 -1760 2100
rect -2020 1980 -1760 2020
rect -2020 1900 -1980 1980
rect -1860 1900 -1760 1980
rect -2020 1860 -1760 1900
rect -2020 1780 -1980 1860
rect -1860 1780 -1760 1860
rect 700 1800 1200 2100
rect -2020 1700 -1760 1780
rect 1000 1300 1200 1800
rect -2020 1060 -1760 1140
rect 1000 1100 2400 1300
rect -2020 980 -1980 1060
rect -1860 980 -1760 1060
rect -2020 940 -1760 980
rect -2020 860 -1980 940
rect -1860 860 -1760 940
rect -2020 820 -1760 860
rect -2020 740 -1980 820
rect -1860 740 -1760 820
rect -2020 700 -1760 740
rect 800 700 2400 1100
rect -508 160 -380 632
rect 1700 300 2400 700
rect 1700 100 1800 300
rect 2000 100 2100 300
rect 2300 100 2400 300
rect 4240 200 4660 300
rect 1700 0 2400 100
rect 1700 -200 1800 0
rect 2000 -200 2100 0
rect 2300 -200 2400 0
rect 1700 -300 2400 -200
rect 4080 100 4780 200
rect 4080 -100 4200 100
rect 4400 -100 4500 100
rect 4700 -100 4780 100
rect 4080 -200 4780 -100
rect 4080 -400 4200 -200
rect 4400 -400 4500 -200
rect 4700 -400 4780 -200
rect 4080 -500 4780 -400
rect -2860 -2620 -2440 -2500
rect -2860 -2700 -1000 -2620
rect -2900 -2800 -1000 -2700
rect -2900 -3000 -2700 -2800
rect -2500 -3000 -2400 -2800
rect -2200 -3000 -2100 -2800
rect -1900 -3000 -1800 -2800
rect -1600 -3000 -1500 -2800
rect -1300 -3000 -1000 -2800
rect -2900 -3200 -1000 -3000
<< via2 >>
rect -1980 2020 -1860 2100
rect -1980 1900 -1860 1980
rect -1980 1780 -1860 1860
rect -1980 980 -1860 1060
rect -1980 860 -1860 940
rect -1980 740 -1860 820
rect 1800 100 2000 300
rect 2100 100 2300 300
rect 1800 -200 2000 0
rect 2100 -200 2300 0
rect 4200 -100 4400 100
rect 4500 -100 4700 100
rect 4200 -400 4400 -200
rect 4500 -400 4700 -200
rect -2700 -3000 -2500 -2800
rect -2400 -3000 -2200 -2800
rect -2100 -3000 -1900 -2800
rect -1800 -3000 -1600 -2800
rect -1500 -3000 -1300 -2800
<< metal3 >>
rect 100 2300 1900 2400
rect -2020 2100 -1820 2140
rect -2020 2020 -1980 2100
rect -1860 2020 -1820 2100
rect -2020 1980 -1820 2020
rect 100 2100 1300 2300
rect 1800 2100 1900 2300
rect 100 2000 1900 2100
rect -2020 1900 -1980 1980
rect -1860 1900 -1820 1980
rect -2020 1860 -1820 1900
rect -2020 1780 -1980 1860
rect -1860 1780 -1820 1860
rect -2020 1700 -1820 1780
rect 1200 1800 1300 2000
rect 1800 1800 1900 2000
rect 1200 1700 1900 1800
rect 1200 1500 1300 1700
rect 1800 1500 1900 1700
rect -2020 1060 -1820 1140
rect -2020 980 -1980 1060
rect -1860 980 -1820 1060
rect -2020 940 -1820 980
rect -2020 860 -1980 940
rect -1860 860 -1820 940
rect 1200 900 1900 1500
rect -2020 820 -1820 860
rect -2020 740 -1980 820
rect -1860 740 -1820 820
rect -2020 700 -1820 740
rect 100 500 1900 900
rect 1700 300 2400 400
rect 1700 100 1800 300
rect 2000 100 2100 300
rect 2300 200 2400 300
rect 2300 100 4780 200
rect 1700 0 4200 100
rect 1700 -200 1800 0
rect 2000 -200 2100 0
rect 2300 -100 4200 0
rect 4400 -100 4500 100
rect 4700 -100 4780 100
rect 2300 -200 2400 -100
rect 1700 -300 2400 -200
rect 2600 -300 2700 -100
rect 2900 -300 3000 -100
rect 3200 -200 4780 -100
rect 3200 -300 4200 -200
rect 1700 -400 4200 -300
rect 4400 -400 4500 -200
rect 4700 -400 4780 -200
rect 1700 -500 2500 -400
rect 2200 -600 2500 -500
rect 2700 -600 2800 -400
rect 3000 -500 4780 -400
rect 3000 -600 3400 -500
rect -700 -800 600 -700
rect 2200 -800 3400 -600
rect -700 -1100 -600 -800
rect -300 -900 200 -800
rect -300 -1100 -200 -900
rect -700 -1200 -200 -1100
rect 100 -1100 200 -900
rect 500 -1100 600 -800
rect 100 -1200 600 -1100
rect -700 -1500 -600 -1200
rect -300 -1300 200 -1200
rect -300 -1500 -200 -1300
rect -700 -1600 -200 -1500
rect 100 -1500 200 -1300
rect 500 -1500 600 -1200
rect 100 -1600 600 -1500
rect -700 -1700 600 -1600
rect -600 -2700 500 -1700
rect -2800 -2800 500 -2700
rect -2800 -3000 -2700 -2800
rect -2500 -3000 -2400 -2800
rect -2200 -3000 -2100 -2800
rect -1900 -3000 -1800 -2800
rect -1600 -3000 -1500 -2800
rect -1300 -3000 500 -2800
rect -2800 -3200 500 -3000
<< via3 >>
rect -1980 2020 -1860 2100
rect 1300 2100 1800 2300
rect -1980 1900 -1860 1980
rect -1980 1780 -1860 1860
rect 1300 1800 1800 2000
rect 1300 1500 1800 1700
rect -1980 980 -1860 1060
rect -1980 860 -1860 940
rect -1980 740 -1860 820
rect 2400 -300 2600 -100
rect 2700 -300 2900 -100
rect 3000 -300 3200 -100
rect 2500 -600 2700 -400
rect 2800 -600 3000 -400
rect -600 -1100 -300 -800
rect -200 -1200 100 -900
rect 200 -1100 500 -800
rect -600 -1500 -300 -1200
rect -200 -1600 100 -1300
rect 200 -1500 500 -1200
<< metal4 >>
rect 1200 2580 4520 3340
rect 1200 2300 1900 2580
rect 4100 2500 4500 2580
rect -2020 2100 -1820 2140
rect -2020 2020 -1980 2100
rect -1860 2020 -1820 2100
rect -2020 1980 -1820 2020
rect -2020 1900 -1980 1980
rect -1860 1900 -1820 1980
rect -2020 1860 -1820 1900
rect -2020 1780 -1980 1860
rect -1860 1780 -1820 1860
rect -2020 1400 -1820 1780
rect 1200 2100 1300 2300
rect 1800 2100 1900 2300
rect 1200 2000 1900 2100
rect 1200 1800 1300 2000
rect 1800 1800 1900 2000
rect 1200 1700 1900 1800
rect 1200 1500 1300 1700
rect 1800 1500 1900 1700
rect 1200 1400 1900 1500
rect -6000 1060 -1820 1400
rect -6000 980 -1980 1060
rect -1860 980 -1820 1060
rect -6000 940 -1820 980
rect -6000 860 -1980 940
rect -1860 860 -1820 940
rect -6000 820 -1820 860
rect -6000 740 -1980 820
rect -1860 740 -1820 820
rect -6000 700 -1820 740
rect -6000 200 -2000 700
rect -6000 -400 -5800 200
rect -4800 0 -2000 200
rect -4800 -20 -4400 0
rect -4800 -400 -4600 -20
rect -2700 -260 -2300 0
rect 2300 -100 3300 0
rect -6000 -12100 -4600 -400
rect 2300 -300 2400 -100
rect 2600 -300 2700 -100
rect 2900 -300 3000 -100
rect 3200 -300 3300 -100
rect 2300 -400 3300 -300
rect 2300 -600 2500 -400
rect 2700 -600 2800 -400
rect 3000 -600 3300 -400
rect 2300 -700 3300 -600
rect -700 -800 600 -700
rect -700 -1100 -600 -800
rect -300 -900 200 -800
rect -300 -1100 -200 -900
rect -700 -1200 -200 -1100
rect 100 -1100 200 -900
rect 500 -1100 600 -800
rect 100 -1200 600 -1100
rect -700 -1500 -600 -1200
rect -300 -1300 200 -1200
rect -300 -1500 -200 -1300
rect -700 -1600 -200 -1500
rect 100 -1500 200 -1300
rect 500 -1500 600 -1200
rect 100 -1600 600 -1500
rect -700 -1700 600 -1600
<< via4 >>
rect -5800 -400 -4800 200
rect -600 -1100 -300 -800
rect -200 -1200 100 -900
rect 200 -1100 500 -800
rect -600 -1500 -300 -1200
rect -200 -1600 100 -1300
rect 200 -1500 500 -1200
<< metal5 >>
rect 7640 3440 10240 4440
rect -6000 200 -4600 400
rect -6800 -400 -5800 200
rect -4800 -400 -4600 200
rect -6000 -600 -4600 -400
use CPW_chunk_W3L5  CPW_chunk_W3L5_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1658705077
transform 1 0 -7800 0 1 -800
box 0 -1000 1200 2400
use CPW_chunk_W3L5  CPW_chunk_W3L5_1
timestamp 1658705077
transform 1 0 -9000 0 1 -800
box 0 -1000 1200 2400
use CPW_chunk_W3L5  CPW_chunk_W3L5_2
timestamp 1658705077
transform 1 0 -10200 0 1 -800
box 0 -1000 1200 2400
use CPW_chunk_W3L5  CPW_chunk_W3L5_3
timestamp 1658705077
transform 1 0 -11400 0 1 -800
box 0 -1000 1200 2400
use CPW_chunk_W3L5  CPW_chunk_W3L5_4
timestamp 1658705077
transform 1 0 -12600 0 1 -800
box 0 -1000 1200 2400
use CPW_chunk_W3L5  CPW_chunk_W3L5_5
timestamp 1658705077
transform 1 0 -13800 0 1 -800
box 0 -1000 1200 2400
use captuner_complete_1  captuner_complete_1_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/COMMON
timestamp 1660736647
transform 1 0 6100 0 1 -800
box -3300 1000 -300 3400
use captuner_complete_1  captuner_complete_1_1
timestamp 1660736647
transform -1 0 -4300 0 1 -3600
box -3300 1000 -300 3400
use nfet_3x_2  nfet_3x_2_0
timestamp 1660736647
transform 1 0 -400 0 1 60
box 0 -60 1292 1380
use nfet_3x_2  nfet_3x_2_1
timestamp 1660736647
transform 1 0 -400 0 -1 2780
box 0 -60 1292 1380
use nfet_3x_2  nfet_3x_2_2
timestamp 1660736647
transform -1 0 -488 0 1 60
box 0 -60 1292 1380
use nfet_3x_2  nfet_3x_2_3
timestamp 1660736647
transform -1 0 -488 0 -1 2780
box 0 -60 1292 1380
use sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top_0 ~/openmpw/pdk_1/sky130A/libs.ref/sky130_fd_pr/mag
timestamp 1649977179
transform 1 0 -7340 0 1 1780
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top_1
timestamp 1649977179
transform 1 0 -11960 0 1 1780
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top_2
timestamp 1649977179
transform 1 0 -3400 0 1 -8100
box 0 0 4498 4610
use sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top  sky130_fd_pr__cap_vpp_11p5x11p7_l1m1m2m3_shieldpom4_top_3
timestamp 1649977179
transform 1 0 -3400 0 1 -12900
box 0 0 4498 4610
use square_ind_0p502n_5GHz  square_ind_0p502n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1658699409
transform 1 0 -1100 0 1 -100
box 200 -13600 13200 -300
use square_ind_1p6n_5GHz  square_ind_1p6n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1658697764
transform -1 0 8040 0 -1 4240
box -200 -19200 19800 1400
use square_ind_2p99n_5GHz  square_ind_2p99n_5GHz_0 ~/openmpw/Project-Yatsuhashi-Chip1/mag/IND
timestamp 1658694498
transform 0 1 -7800 -1 0 -4200
box -1000 -23000 23000 1400
<< end >>
